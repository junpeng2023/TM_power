module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net646;
 wire clknet_1_0__leaf_net646;
 wire clknet_1_1__leaf_net646;
 wire clknet_0_net736;
 wire clknet_1_0__leaf_net736;
 wire clknet_1_1__leaf_net736;
 wire clknet_0_net632;
 wire clknet_1_0__leaf_net632;
 wire clknet_1_1__leaf_net632;
 wire clknet_0_net735;
 wire clknet_1_0__leaf_net735;
 wire clknet_1_1__leaf_net735;
 wire clknet_0_net716;
 wire clknet_1_0__leaf_net716;
 wire clknet_1_1__leaf_net716;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net576;
 wire clknet_1_0__leaf_net576;
 wire clknet_1_1__leaf_net576;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net598;
 wire clknet_1_0__leaf_net598;
 wire clknet_1_1__leaf_net598;
 wire clknet_0_net834;
 wire clknet_1_0__leaf_net834;
 wire clknet_1_1__leaf_net834;
 wire clknet_0_net531;
 wire clknet_1_0__leaf_net531;
 wire clknet_1_1__leaf_net531;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net826;
 wire clknet_1_0__leaf_net826;
 wire clknet_1_1__leaf_net826;
 wire clknet_0_net687;
 wire clknet_1_0__leaf_net687;
 wire clknet_1_1__leaf_net687;
 wire clknet_0_net846;
 wire clknet_1_0__leaf_net846;
 wire clknet_1_1__leaf_net846;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net386;
 wire clknet_1_0__leaf_net386;
 wire clknet_1_1__leaf_net386;
 wire clknet_0_net633;
 wire clknet_1_0__leaf_net633;
 wire clknet_1_1__leaf_net633;
 wire clknet_0_net393;
 wire clknet_1_0__leaf_net393;
 wire clknet_1_1__leaf_net393;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net686;
 wire clknet_1_0__leaf_net686;
 wire clknet_1_1__leaf_net686;
 wire clknet_0_net672;
 wire clknet_1_0__leaf_net672;
 wire clknet_1_1__leaf_net672;
 wire clknet_0_net403;
 wire clknet_1_0__leaf_net403;
 wire clknet_1_1__leaf_net403;
 wire clknet_0_net831;
 wire clknet_1_0__leaf_net831;
 wire clknet_1_1__leaf_net831;
 wire clknet_0_net871;
 wire clknet_1_0__leaf_net871;
 wire clknet_1_1__leaf_net871;
 wire clknet_0_net671;
 wire clknet_1_0__leaf_net671;
 wire clknet_1_1__leaf_net671;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net154;
 wire clknet_1_0__leaf_net154;
 wire clknet_1_1__leaf_net154;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net855;
 wire clknet_1_0__leaf_net855;
 wire clknet_1_1__leaf_net855;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net859;
 wire clknet_1_0__leaf_net859;
 wire clknet_1_1__leaf_net859;
 wire clknet_0_net874;
 wire clknet_1_0__leaf_net874;
 wire clknet_1_1__leaf_net874;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net155;
 wire clknet_1_0__leaf_net155;
 wire clknet_1_1__leaf_net155;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net375;
 wire clknet_1_0__leaf_net375;
 wire clknet_1_1__leaf_net375;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;

 sky130_fd_sc_hd__and2_1 c100 (.A(net37),
    .B(net31),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net27),
    .A1(net33),
    .A2(net22),
    .A3(net18),
    .S0(net992),
    .S1(net38),
    .X(net39));
 sky130_fd_sc_hd__and3_1 c102 (.A(net31),
    .B(net34),
    .C(net37),
    .X(net40));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net23),
    .A1(net38),
    .A2(net35),
    .A3(net25),
    .S0(net40),
    .S1(net984),
    .X(net41));
 sky130_fd_sc_hd__sdfrbp_1 c104 (.CLK(clknet_leaf_6_clk),
    .D(net36),
    .RESET_B(net37),
    .SCD(net40),
    .SCE(net31),
    .Q(net43),
    .Q_N(net42));
 sky130_fd_sc_hd__and2_1 c105 (.A(net779),
    .B(net36),
    .X(net44));
 sky130_fd_sc_hd__and2_0 c106 (.A(net31),
    .B(net19),
    .X(net45));
 sky130_fd_sc_hd__and2_1 c107 (.A(net29),
    .B(net30),
    .X(net46));
 sky130_fd_sc_hd__and2_0 c108 (.A(net45),
    .B(net651),
    .X(net47));
 sky130_fd_sc_hd__dfrbp_1 c109 (.CLK(clknet_leaf_7_clk),
    .D(net40),
    .RESET_B(net31),
    .Q(net876),
    .Q_N(net48));
 sky130_fd_sc_hd__dfbbn_1 c110 (.CLK_N(clknet_leaf_8_clk),
    .D(net44),
    .RESET_B(net903),
    .SET_B(net652),
    .Q(net50),
    .Q_N(net49));
 sky130_fd_sc_hd__and2_1 c111 (.A(net36),
    .B(net768),
    .X(net51));
 sky130_fd_sc_hd__and2_1 c112 (.A(net45),
    .B(net29),
    .X(net52));
 sky130_fd_sc_hd__dfrbp_1 c113 (.CLK(clknet_leaf_8_clk),
    .D(net52),
    .RESET_B(net49),
    .Q(net54),
    .Q_N(net53));
 sky130_fd_sc_hd__dfrtn_1 c114 (.CLK_N(clknet_leaf_8_clk),
    .D(net51),
    .RESET_B(net44),
    .Q(net55));
 sky130_fd_sc_hd__sdfbbn_2 c115 (.CLK_N(clknet_leaf_7_clk),
    .D(net51),
    .RESET_B(net19),
    .SCD(net48),
    .SCE(net47),
    .SET_B(net31),
    .Q(net57),
    .Q_N(net56));
 sky130_fd_sc_hd__or4bb_1 c116 (.A(net939),
    .B(net57),
    .C_N(net29),
    .D_N(net53),
    .X(net58));
 sky130_fd_sc_hd__dfbbn_1 c117 (.CLK_N(clknet_leaf_8_clk),
    .D(net57),
    .RESET_B(net52),
    .SET_B(net58),
    .Q(net862),
    .Q_N(net59));
 sky130_fd_sc_hd__and2_0 c118 (.A(net50),
    .B(net57),
    .X(net830));
 sky130_fd_sc_hd__dfbbp_1 c119 (.CLK(clknet_leaf_7_clk),
    .D(net58),
    .RESET_B(net51),
    .SET_B(net44),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__and3_1 c120 (.A(net61),
    .B(net59),
    .C(net56),
    .X(net62));
 sky130_fd_sc_hd__sdfbbn_1 c121 (.CLK_N(clknet_leaf_7_clk),
    .D(net52),
    .RESET_B(net939),
    .SCD(net62),
    .SCE(net57),
    .SET_B(net61),
    .Q(net835),
    .Q_N(net63));
 sky130_fd_sc_hd__and2_1 c122 (.A(net862),
    .B(net33),
    .X(net827));
 sky130_fd_sc_hd__mux4_1 c123 (.A0(net62),
    .A1(net827),
    .A2(net31),
    .A3(net19),
    .S0(net56),
    .S1(net60),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net47),
    .A1(net30),
    .A2(net827),
    .A3(net56),
    .S0(net64),
    .S1(net980),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net64),
    .A1(net827),
    .A2(net56),
    .A3(net31),
    .S0(net903),
    .S1(net978),
    .X(net66));
 sky130_fd_sc_hd__and3_2 c126 (.A(net769),
    .B(net766),
    .C(net768),
    .X(net857));
 sky130_fd_sc_hd__and2_1 c127 (.A(net821),
    .B(net767),
    .X(net67));
 sky130_fd_sc_hd__mux4_2 c128 (.A0(net768),
    .A1(net67),
    .A2(net763),
    .A3(net769),
    .S0(net901),
    .S1(net794),
    .X(net68));
 sky130_fd_sc_hd__and2_4 c129 (.A(net770),
    .B(net761),
    .X(net69));
 sky130_fd_sc_hd__and2_4 c130 (.A(net805),
    .B(net766),
    .X(net70));
 sky130_fd_sc_hd__or4bb_4 c131 (.A(net821),
    .B(net900),
    .C_N(net816),
    .D_N(net767),
    .X(net71));
 sky130_fd_sc_hd__and2_1 c132 (.A(net819),
    .B(net761),
    .X(net72));
 sky130_fd_sc_hd__and2_1 c133 (.A(net71),
    .B(net783),
    .X(net73));
 sky130_fd_sc_hd__and2_0 c134 (.A(net73),
    .B(net901),
    .X(net74));
 sky130_fd_sc_hd__and3_1 c135 (.A(net72),
    .B(net900),
    .C(net765),
    .X(net75));
 sky130_fd_sc_hd__and3_1 c136 (.A(net901),
    .B(net75),
    .C(net71),
    .X(net76));
 sky130_fd_sc_hd__and3_2 c137 (.A(net75),
    .B(net72),
    .C(net69),
    .X(net77));
 sky130_fd_sc_hd__and2_1 c138 (.A(net763),
    .B(net74),
    .X(net78));
 sky130_fd_sc_hd__and3_2 c139 (.A(net783),
    .B(net75),
    .C(net901),
    .X(net79));
 sky130_fd_sc_hd__a2111o_1 c140 (.A1(net72),
    .A2(net79),
    .B1(net900),
    .C1(net78),
    .D1(net901),
    .X(net80));
 sky130_fd_sc_hd__and3_1 c141 (.A(net764),
    .B(net76),
    .C(net69),
    .X(net81));
 sky130_fd_sc_hd__and3_4 c142 (.A(net81),
    .B(net816),
    .C(net820),
    .X(net82));
 sky130_fd_sc_hd__and2_4 c143 (.A(net82),
    .B(net81),
    .X(net83));
 sky130_fd_sc_hd__and3_4 c144 (.A(net77),
    .B(net771),
    .C(net83),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net78),
    .A1(net73),
    .A2(net764),
    .A3(net82),
    .S0(net769),
    .S1(net69),
    .X(net85));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net80),
    .A1(net85),
    .A2(net83),
    .A3(net72),
    .S0(net73),
    .S1(net82),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c147 (.A(net786),
    .B(net791),
    .C(net771),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c148 (.A(net78),
    .B(net782),
    .X(net88));
 sky130_fd_sc_hd__and3_4 c149 (.A(net767),
    .B(net84),
    .C(net760),
    .X(net89));
 sky130_fd_sc_hd__and2_1 c150 (.A(net791),
    .B(net767),
    .X(net90));
 sky130_fd_sc_hd__and3_1 c151 (.A(net88),
    .B(net768),
    .C(net89),
    .X(net91));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net87),
    .A1(net89),
    .A2(net767),
    .A3(net69),
    .S0(net768),
    .S1(net792),
    .X(net92));
 sky130_fd_sc_hd__and3_1 c153 (.A(net90),
    .B(net87),
    .C(net89),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c154 (.A(net796),
    .B(net68),
    .X(net94));
 sky130_fd_sc_hd__or4bb_2 c155 (.A(net68),
    .B(net90),
    .C_N(net88),
    .D_N(net782),
    .X(net95));
 sky130_fd_sc_hd__a2111o_1 c156 (.A1(net88),
    .A2(net79),
    .B1(net820),
    .C1(net775),
    .D1(net785),
    .X(net96));
 sky130_fd_sc_hd__and2_1 c157 (.A(net788),
    .B(net93),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c158 (.A0(net93),
    .A1(net91),
    .A2(net68),
    .A3(net87),
    .S0(net789),
    .S1(net97),
    .X(net98));
 sky130_fd_sc_hd__a2111o_1 c159 (.A1(net784),
    .A2(net787),
    .B1(net792),
    .C1(net780),
    .D1(net97),
    .X(net99));
 sky130_fd_sc_hd__or4bb_2 c160 (.A(net94),
    .B(net83),
    .C_N(net782),
    .D_N(net787),
    .X(net100));
 sky130_fd_sc_hd__or4bb_4 c161 (.A(net790),
    .B(net792),
    .C_N(net92),
    .D_N(net100),
    .X(net101));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net96),
    .A1(net101),
    .A2(net89),
    .A3(net87),
    .S0(net83),
    .S1(net99),
    .X(net102));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net778),
    .A1(net93),
    .A2(net99),
    .A3(net89),
    .S0(net98),
    .S1(net791),
    .X(net103));
 sky130_fd_sc_hd__a2111o_1 c164 (.A1(net89),
    .A2(net101),
    .B1(net96),
    .C1(net885),
    .D1(net779),
    .X(net104));
 sky130_fd_sc_hd__a2111o_2 c165 (.A1(net95),
    .A2(net791),
    .B1(net97),
    .C1(net104),
    .D1(net79),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net927),
    .A1(net105),
    .A2(net104),
    .A3(net90),
    .S0(net88),
    .S1(net103),
    .X(net106));
 sky130_fd_sc_hd__sdfbbp_1 c167 (.CLK(clknet_leaf_42_clk),
    .D(net100),
    .RESET_B(net106),
    .SCD(net99),
    .SCE(net782),
    .SET_B(net885),
    .Q(net108),
    .Q_N(net107));
 sky130_fd_sc_hd__and3_1 c168 (.A(net771),
    .B(net79),
    .C(net0),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c169 (.A(net91),
    .B(net782),
    .X(net110));
 sky130_fd_sc_hd__and3_2 c170 (.A(net809),
    .B(net79),
    .C(net782),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c171 (.A(net799),
    .B(net109),
    .C(net903),
    .X(net112));
 sky130_fd_sc_hd__and2_0 c172 (.A(net109),
    .B(net903),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c173 (.A(net781),
    .B(net885),
    .C(net107),
    .X(net114));
 sky130_fd_sc_hd__and3_1 c174 (.A(net112),
    .B(net114),
    .C(net900),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c175 (.A(net777),
    .B(net111),
    .C(net112),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c176 (.A(net99),
    .B(net114),
    .C(net110),
    .X(net117));
 sky130_fd_sc_hd__and3_1 c177 (.A(net116),
    .B(net903),
    .C(net782),
    .X(net118));
 sky130_fd_sc_hd__and2_1 c178 (.A(net118),
    .B(net115),
    .X(net119));
 sky130_fd_sc_hd__sdfxbp_1 c179 (.CLK(clknet_leaf_43_clk),
    .D(net110),
    .SCD(net115),
    .SCE(net119),
    .Q(net121),
    .Q_N(net120));
 sky130_fd_sc_hd__and3_2 c180 (.A(net117),
    .B(net118),
    .C(net113),
    .X(net122));
 sky130_fd_sc_hd__sdfxbp_1 c181 (.CLK(clknet_leaf_42_clk),
    .D(net119),
    .SCD(net110),
    .SCE(net111),
    .Q(net123));
 sky130_fd_sc_hd__sdfxtp_1 c182 (.CLK(clknet_leaf_42_clk),
    .D(net946),
    .SCD(net119),
    .SCE(net776),
    .Q(net124));
 sky130_fd_sc_hd__sdfxtp_1 c183 (.CLK(clknet_leaf_43_clk),
    .D(net113),
    .SCD(net122),
    .SCE(net944),
    .Q(net125));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net944),
    .A1(net885),
    .A2(net118),
    .A3(net812),
    .S0(net109),
    .S1(net122),
    .X(net126));
 sky130_fd_sc_hd__sdfxtp_1 c185 (.CLK(clknet_leaf_42_clk),
    .D(net111),
    .SCD(net122),
    .SCE(net115),
    .Q(net127));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(net97),
    .A1(net112),
    .A2(net760),
    .A3(net927),
    .S0(net118),
    .S1(net894),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net79),
    .A1(net109),
    .A2(net112),
    .A3(net900),
    .S0(net122),
    .S1(net894),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net128),
    .A1(net127),
    .A2(net797),
    .A3(net782),
    .S0(net894),
    .S1(clknet_1_0__leaf_net859),
    .X(net130));
 sky130_fd_sc_hd__sdfbbn_1 c189 (.CLK_N(clknet_leaf_5_clk),
    .D(net125),
    .RESET_B(net17),
    .SCD(net77),
    .SCE(net891),
    .SET_B(net122),
    .Q(net131));
 sky130_fd_sc_hd__and3_1 c190 (.A(net1),
    .B(net108),
    .C(net13),
    .X(net132));
 sky130_fd_sc_hd__and3_1 c191 (.A(net818),
    .B(net77),
    .C(net808),
    .X(net133));
 sky130_fd_sc_hd__and3_1 c192 (.A(net90),
    .B(net901),
    .C(net104),
    .X(net134));
 sky130_fd_sc_hd__and3_2 c193 (.A(net131),
    .B(net17),
    .C(net21),
    .X(net135));
 sky130_fd_sc_hd__and3_1 c194 (.A(net18),
    .B(net21),
    .C(net792),
    .X(net136));
 sky130_fd_sc_hd__and2_0 c195 (.A(net134),
    .B(net136),
    .X(net137));
 sky130_fd_sc_hd__and3_2 c196 (.A(net104),
    .B(net812),
    .C(net135),
    .X(net138));
 sky130_fd_sc_hd__and3_1 c197 (.A(net17),
    .B(net804),
    .C(net882),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c198 (.A(net808),
    .B(net108),
    .C(net894),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net20),
    .A1(net804),
    .A2(net21),
    .A3(net12),
    .S0(net135),
    .S1(net892),
    .X(net141));
 sky130_fd_sc_hd__sdfbbn_2 c200 (.CLK_N(clknet_leaf_5_clk),
    .D(net137),
    .RESET_B(net134),
    .SCD(net1),
    .SCE(net125),
    .SET_B(net892),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__sdfbbp_1 c201 (.CLK(clknet_leaf_4_clk),
    .D(net139),
    .RESET_B(net760),
    .SCD(net892),
    .SCE(net141),
    .SET_B(net6),
    .Q(net145),
    .Q_N(net144));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(net782),
    .A1(net787),
    .A2(net122),
    .A3(net895),
    .S0(net882),
    .S1(net142),
    .X(net146));
 sky130_fd_sc_hd__sdfbbn_1 c203 (.CLK_N(clknet_leaf_4_clk),
    .D(net115),
    .RESET_B(net6),
    .SCD(net892),
    .SCE(net143),
    .SET_B(net122),
    .Q(net148),
    .Q_N(net147));
 sky130_fd_sc_hd__or4bb_2 c204 (.A(net812),
    .B(net148),
    .C_N(net142),
    .D_N(net892),
    .X(net149));
 sky130_fd_sc_hd__dfbbn_1 c205 (.CLK_N(clknet_leaf_4_clk),
    .D(net149),
    .RESET_B(net139),
    .SET_B(net976),
    .Q(net151),
    .Q_N(net150));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net148),
    .A1(net143),
    .A2(net892),
    .A3(net882),
    .S0(net139),
    .S1(net808),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net122),
    .A1(net895),
    .A2(net145),
    .A3(net137),
    .S0(net148),
    .S1(clknet_1_0__leaf_net655),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net133),
    .A1(net132),
    .A2(net147),
    .A3(clknet_1_0__leaf_net654),
    .S0(clknet_1_0__leaf_net655),
    .S1(net657),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net6),
    .A1(net892),
    .A2(net121),
    .A3(net147),
    .S0(clknet_1_0__leaf_net859),
    .S1(net656),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c210 (.A(net820),
    .B(net34),
    .C(clknet_1_0__leaf_net859),
    .X(net156));
 sky130_fd_sc_hd__and2_1 c211 (.A(net34),
    .B(net11),
    .X(net157));
 sky130_fd_sc_hd__dfbbn_1 c212 (.CLK_N(clknet_leaf_7_clk),
    .D(net38),
    .RESET_B(net149),
    .SET_B(net652),
    .Q(net159),
    .Q_N(net158));
 sky130_fd_sc_hd__and3_1 c213 (.A(net141),
    .B(net159),
    .C(net928),
    .X(net160));
 sky130_fd_sc_hd__or4bb_2 c214 (.A(net797),
    .B(net903),
    .C_N(net142),
    .D_N(net905),
    .X(net161));
 sky130_fd_sc_hd__and2_1 c215 (.A(net929),
    .B(net12),
    .X(net162));
 sky130_fd_sc_hd__dfbbp_1 c216 (.CLK(clknet_leaf_6_clk),
    .D(clknet_1_1__leaf_net156),
    .RESET_B(net161),
    .SET_B(net940),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__sdfrbp_1 c217 (.CLK(clknet_leaf_6_clk),
    .D(clknet_1_0__leaf_net156),
    .RESET_B(net934),
    .SCD(net928),
    .SCE(net161),
    .Q(net166),
    .Q_N(net165));
 sky130_fd_sc_hd__or4bb_2 c218 (.A(net143),
    .B(net18),
    .C_N(net111),
    .D_N(net160),
    .X(net167));
 sky130_fd_sc_hd__sdfxbp_1 c219 (.CLK(clknet_leaf_6_clk),
    .D(net167),
    .SCD(net18),
    .SCE(net161),
    .Q(net852),
    .Q_N(net168));
 sky130_fd_sc_hd__mux4_2 c220 (.A0(net134),
    .A1(net35),
    .A2(net928),
    .A3(net142),
    .S0(net43),
    .S1(net161),
    .X(net169));
 sky130_fd_sc_hd__sdfxbp_1 c221 (.CLK(clknet_leaf_6_clk),
    .D(net949),
    .SCD(net169),
    .SCE(net162),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__a2111o_1 c222 (.A1(net162),
    .A2(net760),
    .B1(net820),
    .C1(net170),
    .D1(net168),
    .X(net172));
 sky130_fd_sc_hd__sdfxtp_1 c223 (.CLK(clknet_leaf_6_clk),
    .D(net947),
    .SCD(net172),
    .SCE(net169),
    .Q(net173));
 sky130_fd_sc_hd__and2_1 c224 (.A(net161),
    .B(net140),
    .X(net174));
 sky130_fd_sc_hd__and3_1 c225 (.A(net172),
    .B(net174),
    .C(net143),
    .X(net175));
 sky130_fd_sc_hd__and3_2 c226 (.A(net173),
    .B(net165),
    .C(net144),
    .X(net850));
 sky130_fd_sc_hd__and3_1 c227 (.A(net11),
    .B(net173),
    .C(net850),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net43),
    .A1(net149),
    .A2(net174),
    .A3(net850),
    .S0(net175),
    .S1(net176),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net174),
    .A1(net167),
    .A2(net175),
    .A3(net158),
    .S0(net7),
    .S1(net659),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net176),
    .A1(net850),
    .A2(net787),
    .A3(net28),
    .S0(net175),
    .S1(net869),
    .X(net179));
 sky130_fd_sc_hd__and3_1 c231 (.A(net892),
    .B(net54),
    .C(net652),
    .X(net853));
 sky130_fd_sc_hd__or4bb_1 c232 (.A(net787),
    .B(net768),
    .C_N(net57),
    .D_N(clknet_1_1__leaf_net859),
    .X(net180));
 sky130_fd_sc_hd__a2111o_1 c233 (.A1(net159),
    .A2(net63),
    .B1(net807),
    .C1(net56),
    .D1(net853),
    .X(net181));
 sky130_fd_sc_hd__and3_1 c234 (.A(net145),
    .B(net789),
    .C(net22),
    .X(net182));
 sky130_fd_sc_hd__a2111o_1 c235 (.A1(net760),
    .A2(net182),
    .B1(net158),
    .C1(net892),
    .D1(net652),
    .X(net183));
 sky130_fd_sc_hd__and3_1 c236 (.A(net182),
    .B(net853),
    .C(net901),
    .X(net184));
 sky130_fd_sc_hd__or4bb_4 c237 (.A(net183),
    .B(net876),
    .C_N(net768),
    .D_N(net182),
    .X(net185));
 sky130_fd_sc_hd__sdfxtp_1 c238 (.CLK(clknet_leaf_6_clk),
    .D(net157),
    .SCD(net185),
    .SCE(net787),
    .Q(net186));
 sky130_fd_sc_hd__a2111o_1 c239 (.A1(net768),
    .A2(net22),
    .B1(net182),
    .C1(net56),
    .D1(net186),
    .X(net187));
 sky130_fd_sc_hd__sdfbbn_1 c240 (.CLK_N(clknet_leaf_8_clk),
    .D(net46),
    .RESET_B(net145),
    .SCD(net183),
    .SCE(net185),
    .SET_B(net660),
    .Q(net841),
    .Q_N(net188));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net181),
    .A1(net187),
    .A2(net183),
    .A3(net188),
    .S0(net167),
    .S1(net185),
    .X(net189));
 sky130_fd_sc_hd__sdfbbp_1 c242 (.CLK(clknet_leaf_9_clk),
    .D(net184),
    .RESET_B(net46),
    .SCD(net182),
    .SCE(net807),
    .SET_B(net892),
    .Q(net863));
 sky130_fd_sc_hd__and3_1 c243 (.A(net185),
    .B(net187),
    .C(net163),
    .X(net190));
 sky130_fd_sc_hd__mux4_1 c244 (.A0(net180),
    .A1(net185),
    .A2(net168),
    .A3(net182),
    .S0(net59),
    .S1(clknet_1_1__leaf_net859),
    .X(net874));
 sky130_fd_sc_hd__sdfbbn_1 c245 (.CLK_N(clknet_leaf_9_clk),
    .D(net22),
    .RESET_B(clknet_1_0__leaf_net874),
    .SCD(net190),
    .SCE(net167),
    .SET_B(net660),
    .Q(net192),
    .Q_N(net191));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net54),
    .A1(net192),
    .A2(net187),
    .A3(net853),
    .S0(net188),
    .S1(net869),
    .X(net193));
 sky130_fd_sc_hd__mux4_2 c247 (.A0(net164),
    .A1(net193),
    .A2(net852),
    .A3(net190),
    .S0(net22),
    .S1(net185),
    .X(net833));
 sky130_fd_sc_hd__sdfbbn_1 c248 (.CLK_N(clknet_leaf_9_clk),
    .D(net965),
    .RESET_B(net193),
    .SCD(net144),
    .SCE(net157),
    .SET_B(net833),
    .Q(net195),
    .Q_N(net194));
 sky130_fd_sc_hd__a2111o_1 c249 (.A1(net195),
    .A2(net164),
    .B1(clknet_1_0__leaf_net874),
    .C1(net190),
    .D1(net185),
    .X(net196));
 sky130_fd_sc_hd__or4bb_1 c250 (.A(net187),
    .B(net190),
    .C_N(net191),
    .D_N(net194),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net175),
    .A1(clknet_1_0__leaf_net196),
    .A2(net195),
    .A3(net833),
    .S0(net188),
    .S1(net867),
    .X(net197));
 sky130_fd_sc_hd__and2_2 c252 (.A(net769),
    .B(net773),
    .X(net198));
 sky130_fd_sc_hd__and2_4 c253 (.A(net86),
    .B(net74),
    .X(net199));
 sky130_fd_sc_hd__and2_1 c254 (.A(net888),
    .B(net900),
    .X(net200));
 sky130_fd_sc_hd__and2_1 c255 (.A(net76),
    .B(net816),
    .X(net201));
 sky130_fd_sc_hd__and2_4 c256 (.A(net888),
    .B(net86),
    .X(net202));
 sky130_fd_sc_hd__and2_4 c257 (.A(net200),
    .B(net202),
    .X(net203));
 sky130_fd_sc_hd__and3_1 c258 (.A(net816),
    .B(net200),
    .C(net203),
    .X(net204));
 sky130_fd_sc_hd__and3_1 c259 (.A(net201),
    .B(net204),
    .C(net202),
    .X(net205));
 sky130_fd_sc_hd__or4bb_4 c260 (.A(net74),
    .B(net203),
    .C_N(net769),
    .D_N(net202),
    .X(net206));
 sky130_fd_sc_hd__and2_2 c261 (.A(net773),
    .B(net67),
    .X(net207));
 sky130_fd_sc_hd__and3_1 c262 (.A(net766),
    .B(net207),
    .C(net204),
    .X(net208));
 sky130_fd_sc_hd__a2111o_1 c263 (.A1(net203),
    .A2(net201),
    .B1(net888),
    .C1(net76),
    .D1(net86),
    .X(net209));
 sky130_fd_sc_hd__and2_1 c264 (.A(net794),
    .B(net205),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c265 (.A0(net204),
    .A1(net86),
    .A2(net209),
    .A3(net819),
    .S0(net208),
    .S1(net203),
    .X(net211));
 sky130_fd_sc_hd__and3_1 c266 (.A(net210),
    .B(net80),
    .C(net207),
    .X(net212));
 sky130_fd_sc_hd__and3_1 c267 (.A(net207),
    .B(net200),
    .C(net204),
    .X(net213));
 sky130_fd_sc_hd__mux4_2 c268 (.A0(net209),
    .A1(net201),
    .A2(net212),
    .A3(net206),
    .S0(net207),
    .S1(net888),
    .X(net214));
 sky130_fd_sc_hd__sdfxtp_2 c269 (.CLK(clknet_leaf_40_clk),
    .D(net208),
    .SCD(net201),
    .SCE(net214),
    .Q(net215));
 sky130_fd_sc_hd__and3_1 c270 (.A(net67),
    .B(net213),
    .C(net883),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c271 (.A0(net216),
    .A1(net932),
    .A2(net213),
    .A3(net201),
    .S0(net83),
    .S1(net207),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(net205),
    .A1(net907),
    .A2(net771),
    .A3(net214),
    .S0(net204),
    .S1(net883),
    .X(net218));
 sky130_fd_sc_hd__and2_1 c273 (.A(net204),
    .B(net888),
    .X(net219));
 sky130_fd_sc_hd__and2_1 c274 (.A(net771),
    .B(net885),
    .X(net220));
 sky130_fd_sc_hd__and2_1 c275 (.A(net94),
    .B(net100),
    .X(net221));
 sky130_fd_sc_hd__and2_1 c276 (.A(net775),
    .B(net780),
    .X(net222));
 sky130_fd_sc_hd__and2_1 c277 (.A(net220),
    .B(net219),
    .X(net223));
 sky130_fd_sc_hd__and2_4 c278 (.A(net203),
    .B(net81),
    .X(net224));
 sky130_fd_sc_hd__and2_1 c279 (.A(net96),
    .B(net101),
    .X(net225));
 sky130_fd_sc_hd__mux4_2 c280 (.A0(net212),
    .A1(net204),
    .A2(net108),
    .A3(net202),
    .S0(net219),
    .S1(net220),
    .X(net226));
 sky130_fd_sc_hd__dfrtp_4 c281 (.CLK(clknet_leaf_41_clk),
    .D(net222),
    .RESET_B(net226),
    .Q(net227));
 sky130_fd_sc_hd__and3_4 c282 (.A(net200),
    .B(net212),
    .C(net220),
    .X(net228));
 sky130_fd_sc_hd__dfbbn_1 c283 (.CLK_N(clknet_leaf_41_clk),
    .D(net106),
    .RESET_B(net98),
    .SET_B(net226),
    .Q(net230),
    .Q_N(net229));
 sky130_fd_sc_hd__and2_1 c284 (.A(net223),
    .B(net792),
    .X(net231));
 sky130_fd_sc_hd__and3_2 c285 (.A(net222),
    .B(net96),
    .C(net224),
    .X(net232));
 sky130_fd_sc_hd__and3_4 c286 (.A(net219),
    .B(net223),
    .C(net229),
    .X(net233));
 sky130_fd_sc_hd__dfrtp_4 c287 (.CLK(clknet_leaf_37_clk),
    .D(net231),
    .RESET_B(net232),
    .Q(net234));
 sky130_fd_sc_hd__sdfbbp_1 c288 (.CLK(clknet_leaf_40_clk),
    .D(net226),
    .RESET_B(net228),
    .SCD(net223),
    .SCE(net198),
    .SET_B(net888),
    .Q(net236),
    .Q_N(net235));
 sky130_fd_sc_hd__and2_0 c289 (.A(net234),
    .B(net235),
    .X(net237));
 sky130_fd_sc_hd__a2111o_4 c290 (.A1(net236),
    .A2(net219),
    .B1(net232),
    .C1(net221),
    .D1(net883),
    .X(net825));
 sky130_fd_sc_hd__sdfbbn_2 c291 (.CLK_N(clknet_leaf_0_clk),
    .D(net227),
    .RESET_B(net233),
    .SCD(net226),
    .SCE(net237),
    .SET_B(net825),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net237),
    .A1(net239),
    .A2(net775),
    .A3(net234),
    .S0(net225),
    .S1(net779),
    .X(net240));
 sky130_fd_sc_hd__mux4_2 c293 (.A0(net225),
    .A1(net816),
    .A2(net220),
    .A3(net240),
    .S0(net222),
    .S1(net238),
    .X(net832));
 sky130_fd_sc_hd__and2_1 c294 (.A(net240),
    .B(net770),
    .X(net241));
 sky130_fd_sc_hd__dfbbn_1 c295 (.CLK_N(clknet_leaf_0_clk),
    .D(net241),
    .RESET_B(net228),
    .SET_B(net888),
    .Q(net242));
 sky130_fd_sc_hd__and3_1 c296 (.A(net774),
    .B(net103),
    .C(net883),
    .X(net243));
 sky130_fd_sc_hd__and2_1 c297 (.A(net114),
    .B(net112),
    .X(net244));
 sky130_fd_sc_hd__and3_1 c298 (.A(net221),
    .B(net779),
    .C(net883),
    .X(net245));
 sky130_fd_sc_hd__a2111o_1 c299 (.A1(net242),
    .A2(net243),
    .B1(net789),
    .C1(net234),
    .D1(net241),
    .X(net246));
 sky130_fd_sc_hd__sdfbbn_1 c300 (.CLK_N(clknet_leaf_43_clk),
    .D(net243),
    .RESET_B(net246),
    .SCD(net120),
    .SCE(net908),
    .SET_B(net234),
    .Q(net247));
 sky130_fd_sc_hd__dfbbp_1 c301 (.CLK(clknet_leaf_0_clk),
    .D(net246),
    .RESET_B(net103),
    .SET_B(net832),
    .Q(net248));
 sky130_fd_sc_hd__and3_2 c302 (.A(net245),
    .B(net114),
    .C(net103),
    .X(net249));
 sky130_fd_sc_hd__and2_0 c303 (.A(net776),
    .B(net221),
    .X(net250));
 sky130_fd_sc_hd__and3_1 c304 (.A(net247),
    .B(net244),
    .C(net771),
    .X(net251));
 sky130_fd_sc_hd__sdfxbp_1 c305 (.CLK(clknet_leaf_0_clk),
    .D(net103),
    .SCD(net249),
    .SCE(net238),
    .Q(net252));
 sky130_fd_sc_hd__sdfxbp_1 c306 (.CLK(clknet_leaf_1_clk),
    .D(net251),
    .SCD(net249),
    .SCE(net932),
    .Q(net254),
    .Q_N(net253));
 sky130_fd_sc_hd__sdfbbp_1 c307 (.CLK(clknet_leaf_0_clk),
    .D(net250),
    .RESET_B(net251),
    .SCD(net241),
    .SCE(net888),
    .SET_B(net112),
    .Q(net256),
    .Q_N(net255));
 sky130_fd_sc_hd__a2111o_1 c308 (.A1(net93),
    .A2(net800),
    .B1(net224),
    .C1(net77),
    .D1(net888),
    .X(net257));
 sky130_fd_sc_hd__sdfbbn_1 c309 (.CLK_N(clknet_leaf_0_clk),
    .D(net252),
    .RESET_B(net251),
    .SCD(net257),
    .SCE(net244),
    .SET_B(net241),
    .Q(net258));
 sky130_fd_sc_hd__sdfbbn_1 c310 (.CLK_N(clknet_leaf_0_clk),
    .D(net256),
    .RESET_B(net832),
    .SCD(net244),
    .SCE(net246),
    .SET_B(clknet_1_0__leaf_net859),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(net248),
    .A1(net100),
    .A2(net259),
    .A3(net249),
    .S0(net246),
    .S1(net257),
    .X(net261));
 sky130_fd_sc_hd__sdfbbp_1 c312 (.CLK(clknet_leaf_0_clk),
    .D(net257),
    .RESET_B(clknet_1_0__leaf_net130),
    .SCD(net249),
    .SCE(net103),
    .SET_B(net663),
    .Q(net263),
    .Q_N(net262));
 sky130_fd_sc_hd__and3_1 c313 (.A(net258),
    .B(net260),
    .C(net257),
    .X(net264));
 sky130_fd_sc_hd__mux4_2 c314 (.A0(net257),
    .A1(net264),
    .A2(net259),
    .A3(net215),
    .S0(net262),
    .S1(net985),
    .X(net265));
 sky130_fd_sc_hd__and3_1 c315 (.A(net244),
    .B(net803),
    .C(net135),
    .X(net266));
 sky130_fd_sc_hd__sdfxtp_1 c316 (.CLK(clknet_leaf_3_clk),
    .D(clknet_1_1__leaf_net155),
    .SCD(net13),
    .SCE(net233),
    .Q(net267));
 sky130_fd_sc_hd__and3_2 c317 (.A(net936),
    .B(net243),
    .C(net207),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net268),
    .A1(net239),
    .A2(net825),
    .A3(net253),
    .S0(clknet_1_0__leaf_net654),
    .S1(clknet_1_0__leaf_net655),
    .X(net269));
 sky130_fd_sc_hd__sdfxtp_1 c319 (.CLK(clknet_leaf_43_clk),
    .D(net268),
    .SCD(net77),
    .SCE(net888),
    .Q(net270));
 sky130_fd_sc_hd__and3_1 c320 (.A(net267),
    .B(net903),
    .C(net657),
    .X(net271));
 sky130_fd_sc_hd__sdfrtn_1 c321 (.CLK_N(clknet_leaf_4_clk),
    .D(net271),
    .RESET_B(net268),
    .SCD(net906),
    .SCE(net804),
    .Q(net272));
 sky130_fd_sc_hd__and3_1 c322 (.A(net199),
    .B(net272),
    .C(net120),
    .X(net273));
 sky130_fd_sc_hd__and3_2 c323 (.A(net273),
    .B(net215),
    .C(net238),
    .X(net274));
 sky130_fd_sc_hd__sdfxtp_1 c324 (.CLK(clknet_leaf_43_clk),
    .D(net272),
    .SCD(net244),
    .SCE(net268),
    .Q(net845));
 sky130_fd_sc_hd__a2111o_1 c325 (.A1(net896),
    .A2(clknet_1_0__leaf_net154),
    .B1(net274),
    .C1(net883),
    .D1(net77),
    .X(net275));
 sky130_fd_sc_hd__a2111o_1 c326 (.A1(net273),
    .A2(net271),
    .B1(net901),
    .C1(net272),
    .D1(net896),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c327 (.A(net270),
    .B(net207),
    .C(net271),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net804),
    .A1(net249),
    .A2(net273),
    .A3(clknet_1_0__leaf_net275),
    .S0(net896),
    .S1(net277),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net277),
    .A1(clknet_1_1__leaf_net275),
    .A2(net265),
    .A3(clknet_1_0__leaf_net155),
    .S0(net664),
    .S1(net666),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(clknet_1_0__leaf_net275),
    .A1(net761),
    .A2(net273),
    .A3(net239),
    .S0(net896),
    .S1(net656),
    .X(net280));
 sky130_fd_sc_hd__a2111o_1 c331 (.A1(clknet_1_1__leaf_net275),
    .A2(net896),
    .B1(net7),
    .C1(net665),
    .D1(net667),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net274),
    .A1(net243),
    .A2(net21),
    .A3(net896),
    .S0(net664),
    .S1(net666),
    .X(net282));
 sky130_fd_sc_hd__sdfrtp_1 c333 (.CLK(clknet_leaf_2_clk),
    .D(net282),
    .RESET_B(net272),
    .SCD(net896),
    .SCE(net983),
    .Q(net283));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(clknet_1_1__leaf_net280),
    .A1(net268),
    .A2(net271),
    .A3(net274),
    .S0(net896),
    .S1(net657),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_0__leaf_net280),
    .A1(net283),
    .A2(net802),
    .A3(net265),
    .S0(net228),
    .S1(clknet_1_1__leaf_net275),
    .X(net285));
 sky130_fd_sc_hd__and3_1 c336 (.A(net239),
    .B(net276),
    .C(net875),
    .X(net286));
 sky130_fd_sc_hd__and3_2 c337 (.A(net35),
    .B(net107),
    .C(net896),
    .X(net287));
 sky130_fd_sc_hd__and3_1 c338 (.A(net132),
    .B(net286),
    .C(net896),
    .X(net288));
 sky130_fd_sc_hd__and3_2 c339 (.A(net276),
    .B(net7),
    .C(net891),
    .X(net289));
 sky130_fd_sc_hd__and3_1 c340 (.A(net160),
    .B(net897),
    .C(net163),
    .X(net290));
 sky130_fd_sc_hd__and2_1 c341 (.A(net207),
    .B(net287),
    .X(net291));
 sky130_fd_sc_hd__dfbbn_1 c342 (.CLK_N(clknet_leaf_13_clk),
    .D(net254),
    .RESET_B(net290),
    .SET_B(net891),
    .Q(net293),
    .Q_N(net292));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net135),
    .A1(net27),
    .A2(net224),
    .A3(net290),
    .S0(net7),
    .S1(net897),
    .X(net294));
 sky130_fd_sc_hd__and3_1 c344 (.A(net293),
    .B(net289),
    .C(net899),
    .X(net872));
 sky130_fd_sc_hd__and3_1 c345 (.A(net286),
    .B(net135),
    .C(net289),
    .X(net295));
 sky130_fd_sc_hd__dfbbn_1 c346 (.CLK_N(clknet_leaf_3_clk),
    .D(net7),
    .RESET_B(net291),
    .SET_B(net290),
    .Q(net297),
    .Q_N(net296));
 sky130_fd_sc_hd__mux4_2 c347 (.A0(net108),
    .A1(net903),
    .A2(net27),
    .A3(net882),
    .S0(net287),
    .S1(net670),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net288),
    .A1(net174),
    .A2(net132),
    .A3(net897),
    .S0(net27),
    .S1(clknet_1_0__leaf_net655),
    .X(net299));
 sky130_fd_sc_hd__and2_1 c349 (.A(net803),
    .B(net832),
    .X(net300));
 sky130_fd_sc_hd__and3_1 c350 (.A(net295),
    .B(net872),
    .C(net660),
    .X(net838));
 sky130_fd_sc_hd__and3_1 c351 (.A(net838),
    .B(net803),
    .C(net670),
    .X(net301));
 sky130_fd_sc_hd__or4bb_4 c352 (.A(net121),
    .B(net897),
    .C_N(net286),
    .D_N(net107),
    .X(net822));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net301),
    .A1(net287),
    .A2(net838),
    .A3(net292),
    .S0(net882),
    .S1(net670),
    .X(net302));
 sky130_fd_sc_hd__sdfbbn_1 c354 (.CLK_N(clknet_leaf_13_clk),
    .D(net290),
    .RESET_B(net27),
    .SCD(net968),
    .SCE(net897),
    .SET_B(net825),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net304),
    .A1(net301),
    .A2(net822),
    .A3(net289),
    .S0(net238),
    .S1(net658),
    .X(net305));
 sky130_fd_sc_hd__and3_1 c356 (.A(net295),
    .B(net659),
    .C(clknet_1_0__leaf_net672),
    .X(net831));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net789),
    .A1(net822),
    .A2(net833),
    .A3(net838),
    .S0(clknet_1_0__leaf_net831),
    .S1(net867),
    .X(net871));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_0__leaf_net871),
    .A1(clknet_1_1__leaf_net196),
    .A2(net830),
    .A3(net872),
    .S0(net867),
    .S1(net847),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net57),
    .A1(clknet_1_1__leaf_net196),
    .A2(clknet_1_0__leaf_net871),
    .A3(clknet_1_1__leaf_net831),
    .S0(net841),
    .S1(net661),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net193),
    .A1(net167),
    .A2(clknet_1_0__leaf_net871),
    .A3(net899),
    .S0(clknet_1_0__leaf_net196),
    .S1(net847),
    .X(net308));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net186),
    .A1(net164),
    .A2(net841),
    .A3(clknet_1_0__leaf_net871),
    .S0(net853),
    .S1(net673),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net807),
    .A1(net779),
    .A2(clknet_1_0__leaf_net831),
    .A3(net833),
    .S0(net828),
    .S1(net674),
    .X(net861));
 sky130_fd_sc_hd__and2_2 c378 (.A(net80),
    .B(net210),
    .X(net310));
 sky130_fd_sc_hd__a2111o_4 c379 (.A1(net900),
    .A2(net310),
    .B1(net765),
    .C1(net198),
    .D1(net662),
    .X(net311));
 sky130_fd_sc_hd__and2_1 c380 (.A(net75),
    .B(net310),
    .X(net312));
 sky130_fd_sc_hd__and2_2 c381 (.A(net201),
    .B(net83),
    .X(net313));
 sky130_fd_sc_hd__and2_0 c382 (.A(net761),
    .B(net82),
    .X(net314));
 sky130_fd_sc_hd__dfbbp_1 c383 (.CLK(clknet_leaf_39_clk),
    .D(net312),
    .RESET_B(net313),
    .SET_B(net889),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__dfrtp_4 c384 (.CLK(clknet_leaf_39_clk),
    .D(net210),
    .RESET_B(net312),
    .Q(net317));
 sky130_fd_sc_hd__and2_1 c385 (.A(net765),
    .B(net317),
    .X(net318));
 sky130_fd_sc_hd__and2_2 c386 (.A(net310),
    .B(net318),
    .X(net319));
 sky130_fd_sc_hd__and2_1 c387 (.A(net889),
    .B(net215),
    .X(net320));
 sky130_fd_sc_hd__sdfxbp_1 c388 (.CLK(clknet_leaf_39_clk),
    .D(net987),
    .SCD(net319),
    .SCE(net311),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__and2_1 c389 (.A(net313),
    .B(net317),
    .X(net323));
 sky130_fd_sc_hd__sdfrtp_1 c390 (.CLK(clknet_leaf_39_clk),
    .D(net964),
    .RESET_B(net942),
    .SCD(net319),
    .SCE(net889),
    .Q(net324));
 sky130_fd_sc_hd__dfsbp_1 c391 (.CLK(clknet_leaf_39_clk),
    .D(net943),
    .SET_B(net312),
    .Q(net326),
    .Q_N(net325));
 sky130_fd_sc_hd__sdfxbp_1 c392 (.CLK(clknet_leaf_39_clk),
    .D(net987),
    .SCD(net311),
    .SCE(net889),
    .Q(net328),
    .Q_N(net327));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net326),
    .A1(net320),
    .A2(net311),
    .A3(net319),
    .S0(net313),
    .S1(net889),
    .X(net329));
 sky130_fd_sc_hd__and2_0 c394 (.A(net323),
    .B(net327),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net318),
    .A1(net320),
    .A2(net210),
    .A3(net319),
    .S0(net324),
    .S1(net675),
    .X(net331));
 sky130_fd_sc_hd__sdfxtp_1 c396 (.CLK(clknet_leaf_39_clk),
    .D(net311),
    .SCD(net961),
    .SCE(net676),
    .Q(net332));
 sky130_fd_sc_hd__mux4_1 c397 (.A0(net324),
    .A1(net330),
    .A2(net315),
    .A3(net310),
    .S0(net317),
    .S1(net676),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net328),
    .A1(net332),
    .A2(net333),
    .A3(net310),
    .S0(net915),
    .S1(net676),
    .X(net334));
 sky130_fd_sc_hd__and2_1 c399 (.A(net816),
    .B(net310),
    .X(net335));
 sky130_fd_sc_hd__dfsbp_1 c400 (.CLK(clknet_leaf_37_clk),
    .D(net217),
    .SET_B(net313),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__and2_0 c401 (.A(net230),
    .B(net313),
    .X(net338));
 sky130_fd_sc_hd__sdfrtp_4 c402 (.CLK(clknet_leaf_40_clk),
    .D(net335),
    .RESET_B(net83),
    .SCD(net227),
    .SCE(net229),
    .Q(net339));
 sky130_fd_sc_hd__sdfxtp_1 c403 (.CLK(clknet_leaf_38_clk),
    .D(net333),
    .SCD(net230),
    .SCE(net795),
    .Q(net340));
 sky130_fd_sc_hd__mux4_1 c404 (.A0(net780),
    .A1(net912),
    .A2(net231),
    .A3(net69),
    .S0(net215),
    .S1(net313),
    .X(net341));
 sky130_fd_sc_hd__and3_1 c405 (.A(net340),
    .B(net816),
    .C(net678),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c406 (.A0(net335),
    .A1(net232),
    .A2(net340),
    .A3(net101),
    .S0(net336),
    .S1(net678),
    .X(net343));
 sky130_fd_sc_hd__sdfsbp_1 c407 (.CLK(clknet_leaf_38_clk),
    .D(net230),
    .SCD(net982),
    .SCE(net228),
    .SET_B(net933),
    .Q(net345),
    .Q_N(net344));
 sky130_fd_sc_hd__sdfxtp_1 c408 (.CLK(clknet_leaf_38_clk),
    .D(net951),
    .SCD(net335),
    .SCE(net952),
    .Q(net346));
 sky130_fd_sc_hd__and2_1 c409 (.A(net346),
    .B(net337),
    .X(net347));
 sky130_fd_sc_hd__and3_2 c410 (.A(net95),
    .B(net347),
    .C(net901),
    .X(net348));
 sky130_fd_sc_hd__dfstp_1 c411 (.CLK(clknet_leaf_36_clk),
    .D(net231),
    .SET_B(net935),
    .Q(net349));
 sky130_fd_sc_hd__dfstp_1 c412 (.CLK(clknet_leaf_37_clk),
    .D(net948),
    .SET_B(net319),
    .Q(net350));
 sky130_fd_sc_hd__and3_1 c413 (.A(net101),
    .B(net84),
    .C(net349),
    .X(net351));
 sky130_fd_sc_hd__or4bb_1 c414 (.A(net337),
    .B(net101),
    .C_N(net350),
    .D_N(net313),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net352),
    .A1(net339),
    .A2(net348),
    .A3(net340),
    .S0(net347),
    .S1(net889),
    .X(net353));
 sky130_fd_sc_hd__and3_1 c416 (.A(net353),
    .B(net350),
    .C(net352),
    .X(net354));
 sky130_fd_sc_hd__or4bb_2 c417 (.A(net345),
    .B(net354),
    .C_N(net350),
    .D_N(net347),
    .X(net355));
 sky130_fd_sc_hd__and2_2 c418 (.A(net340),
    .B(net677),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net198),
    .A1(net352),
    .A2(net311),
    .A3(net356),
    .S0(net350),
    .S1(net677),
    .X(net357));
 sky130_fd_sc_hd__and2_2 c420 (.A(net98),
    .B(net680),
    .X(net358));
 sky130_fd_sc_hd__and3_1 c421 (.A(net100),
    .B(net215),
    .C(net883),
    .X(net359));
 sky130_fd_sc_hd__and3_2 c422 (.A(net354),
    .B(net359),
    .C(net83),
    .X(net842));
 sky130_fd_sc_hd__sdfsbp_1 c423 (.CLK(clknet_leaf_1_clk),
    .D(net347),
    .SCD(net879),
    .SCE(net224),
    .SET_B(net354),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net351),
    .A1(net265),
    .A2(net311),
    .A3(net251),
    .S0(net879),
    .S1(clknet_1_0__leaf_net859),
    .X(net362));
 sky130_fd_sc_hd__dfbbn_1 c425 (.CLK_N(clknet_leaf_37_clk),
    .D(net224),
    .RESET_B(net228),
    .SET_B(net682),
    .Q(net364),
    .Q_N(net363));
 sky130_fd_sc_hd__sdfbbn_1 c426 (.CLK_N(clknet_leaf_36_clk),
    .D(net811),
    .RESET_B(net955),
    .SCD(net234),
    .SCE(net311),
    .SET_B(net894),
    .Q(net839),
    .Q_N(net365));
 sky130_fd_sc_hd__and3_1 c427 (.A(net358),
    .B(net224),
    .C(net365),
    .X(net366));
 sky130_fd_sc_hd__dfbbn_2 c428 (.CLK_N(clknet_leaf_1_clk),
    .D(net0),
    .RESET_B(net100),
    .SET_B(net311),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__sdfstp_1 c429 (.CLK(clknet_leaf_1_clk),
    .D(net310),
    .SCD(net251),
    .SCE(net802),
    .SET_B(net367),
    .Q(net369));
 sky130_fd_sc_hd__or4bb_4 c430 (.A(net364),
    .B(net234),
    .C_N(net367),
    .D_N(net369),
    .X(net370));
 sky130_fd_sc_hd__a2111o_1 c431 (.A1(net350),
    .A2(net366),
    .B1(net105),
    .C1(net355),
    .D1(net370),
    .X(net371));
 sky130_fd_sc_hd__a2111o_4 c432 (.A1(net366),
    .A2(net370),
    .B1(net368),
    .C1(net358),
    .D1(net811),
    .X(net372));
 sky130_fd_sc_hd__or4bb_4 c433 (.A(net369),
    .B(net347),
    .C_N(net367),
    .D_N(net372),
    .X(net844));
 sky130_fd_sc_hd__a2111o_1 c434 (.A1(net105),
    .A2(net839),
    .B1(net761),
    .C1(net310),
    .D1(clknet_1_1__leaf_net130),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net340),
    .A1(net350),
    .A2(net358),
    .A3(net310),
    .S0(net844),
    .S1(net370),
    .X(net374));
 sky130_fd_sc_hd__a2111o_1 c436 (.A1(net372),
    .A2(net358),
    .B1(net367),
    .C1(clknet_1_0__leaf_net130),
    .D1(net683),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net359),
    .A1(clknet_1_0__leaf_net375),
    .A2(net98),
    .A3(net105),
    .S0(net681),
    .S1(net683),
    .X(net376));
 sky130_fd_sc_hd__sdfstp_2 c438 (.CLK(clknet_leaf_35_clk),
    .D(net368),
    .SCD(clknet_1_1__leaf_net373),
    .SCE(net902),
    .SET_B(net249),
    .Q(net377));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net377),
    .A1(net368),
    .A2(clknet_1_0__leaf_net373),
    .A3(net372),
    .S0(net370),
    .S1(net979),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net844),
    .A1(net377),
    .A2(net310),
    .A3(net679),
    .S0(net684),
    .S1(net945),
    .X(net379));
 sky130_fd_sc_hd__dfbbp_1 c441 (.CLK(clknet_leaf_3_clk),
    .D(net249),
    .RESET_B(net358),
    .SET_B(net265),
    .Q(net381),
    .Q_N(net380));
 sky130_fd_sc_hd__and3_1 c442 (.A(net792),
    .B(net380),
    .C(net668),
    .X(net382));
 sky130_fd_sc_hd__and3_1 c443 (.A(net785),
    .B(net265),
    .C(clknet_1_0__leaf_net655),
    .X(net383));
 sky130_fd_sc_hd__and3_2 c444 (.A(net802),
    .B(net151),
    .C(net761),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net882),
    .A1(net770),
    .A2(net851),
    .A3(net844),
    .S0(net21),
    .S1(net665),
    .X(net384));
 sky130_fd_sc_hd__sdfxbp_1 c446 (.CLK(clknet_leaf_23_clk),
    .D(net902),
    .SCD(clknet_1_1__leaf_net281),
    .SCE(clknet_1_1__leaf_net686),
    .Q(net873),
    .Q_N(net385));
 sky130_fd_sc_hd__and3_1 c447 (.A(net890),
    .B(net274),
    .C(clknet_1_1__leaf_net654),
    .X(net855));
 sky130_fd_sc_hd__or4bb_4 c448 (.A(net885),
    .B(net21),
    .C_N(net898),
    .D_N(clknet_1_0__leaf_net687),
    .X(net386));
 sky130_fd_sc_hd__sdfxbp_1 c449 (.CLK(clknet_leaf_14_clk),
    .D(net381),
    .SCD(clknet_1_0__leaf_net281),
    .SCE(clknet_1_0__leaf_net386),
    .Q(net388),
    .Q_N(net387));
 sky130_fd_sc_hd__or4bb_1 c450 (.A(net370),
    .B(net388),
    .C_N(net901),
    .D_N(clknet_1_0__leaf_net386),
    .X(net389));
 sky130_fd_sc_hd__sdfbbp_1 c451 (.CLK(clknet_leaf_2_clk),
    .D(net266),
    .RESET_B(clknet_1_0__leaf_net386),
    .SCD(net274),
    .SCE(net974),
    .SET_B(net802),
    .Q(net391),
    .Q_N(net390));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(net265),
    .A1(net371),
    .A2(clknet_1_0__leaf_net386),
    .A3(net356),
    .S0(clknet_1_1__leaf_net389),
    .S1(net377),
    .X(net392));
 sky130_fd_sc_hd__a2111o_1 c453 (.A1(net215),
    .A2(net390),
    .B1(clknet_1_0__leaf_net386),
    .C1(net898),
    .D1(net665),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net383),
    .A1(net372),
    .A2(clknet_1_0__leaf_net855),
    .A3(net832),
    .S0(clknet_1_1__leaf_net393),
    .S1(net390),
    .X(net394));
 sky130_fd_sc_hd__a2111o_1 c455 (.A1(net387),
    .A2(clknet_1_1__leaf_net389),
    .B1(clknet_1_1__leaf_net386),
    .C1(net274),
    .D1(net688),
    .X(net826));
 sky130_fd_sc_hd__sdfxtp_1 c456 (.CLK(clknet_leaf_11_clk),
    .D(net382),
    .SCD(clknet_1_1__leaf_net826),
    .SCE(clknet_1_1__leaf_net859),
    .Q(net849));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net361),
    .A1(net851),
    .A2(clknet_1_1__leaf_net389),
    .A3(net387),
    .S0(net668),
    .S1(net689),
    .X(net395));
 sky130_fd_sc_hd__and3_1 c458 (.A(clknet_1_1__leaf_net154),
    .B(clknet_1_0__leaf_net686),
    .C(clknet_1_0__leaf_net687),
    .X(net396));
 sky130_fd_sc_hd__and3_1 c459 (.A(clknet_1_0__leaf_net393),
    .B(net274),
    .C(clknet_1_0__leaf_net386),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net397),
    .A1(net13),
    .A2(net360),
    .A3(net370),
    .S0(net265),
    .S1(net885),
    .X(net398));
 sky130_fd_sc_hd__a2111o_1 c461 (.A1(net396),
    .A2(clknet_1_0__leaf_net855),
    .B1(clknet_1_0__leaf_net386),
    .C1(net898),
    .D1(net894),
    .X(net399));
 sky130_fd_sc_hd__sdfbbn_1 c462 (.CLK_N(clknet_leaf_12_clk),
    .D(net300),
    .RESET_B(net885),
    .SCD(net288),
    .SCE(net28),
    .SET_B(clknet_1_0__leaf_net671),
    .Q(net401),
    .Q_N(net400));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net395),
    .A1(net300),
    .A2(net891),
    .A3(net296),
    .S0(net914),
    .S1(clknet_1_1__leaf_net655),
    .X(net402));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(net293),
    .A1(net289),
    .A2(net851),
    .A3(net28),
    .S0(clknet_1_0__leaf_net671),
    .S1(clknet_1_0__leaf_net672),
    .X(net403));
 sky130_fd_sc_hd__a2111o_1 c465 (.A1(net297),
    .A2(clknet_1_1__leaf_net855),
    .B1(net882),
    .C1(net289),
    .D1(net875),
    .X(net404));
 sky130_fd_sc_hd__a2111o_1 c466 (.A1(net291),
    .A2(net28),
    .B1(clknet_1_0__leaf_net386),
    .C1(net679),
    .D1(clknet_1_1__leaf_net687),
    .X(net846));
 sky130_fd_sc_hd__sdfbbn_1 c467 (.CLK_N(clknet_leaf_14_clk),
    .D(net169),
    .RESET_B(net891),
    .SCD(net902),
    .SCE(clknet_1_0__leaf_net404),
    .SET_B(net12),
    .Q(net405));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net28),
    .A1(net852),
    .A2(net832),
    .A3(net882),
    .S0(clknet_1_1__leaf_net404),
    .S1(net899),
    .X(net406));
 sky130_fd_sc_hd__a2111o_1 c469 (.A1(net883),
    .A2(net913),
    .B1(net851),
    .C1(clknet_1_0__leaf_net386),
    .D1(net694),
    .X(net407));
 sky130_fd_sc_hd__sdfbbp_1 c470 (.CLK(clknet_leaf_13_clk),
    .D(net401),
    .RESET_B(net368),
    .SCD(clknet_1_1__leaf_net404),
    .SCE(net289),
    .SET_B(net938),
    .Q(net409),
    .Q_N(net408));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net289),
    .A1(clknet_1_0__leaf_net846),
    .A2(net300),
    .A3(net885),
    .S0(clknet_1_1__leaf_net671),
    .S1(clknet_1_1__leaf_net687),
    .X(net410));
 sky130_fd_sc_hd__sdfbbn_1 c472 (.CLK_N(clknet_leaf_13_clk),
    .D(clknet_1_0__leaf_net404),
    .RESET_B(net956),
    .SCD(net409),
    .SCE(net224),
    .SET_B(net959),
    .Q(net843));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net388),
    .A1(net300),
    .A2(net408),
    .A3(net291),
    .S0(clknet_1_1__leaf_net859),
    .S1(net848),
    .X(net411));
 sky130_fd_sc_hd__sdfbbn_1 c474 (.CLK_N(clknet_leaf_12_clk),
    .D(net358),
    .RESET_B(clknet_1_1__leaf_net404),
    .SCD(net24),
    .SCE(net899),
    .SET_B(net860),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__a2111o_1 c475 (.A1(net287),
    .A2(net388),
    .B1(clknet_1_0__leaf_net386),
    .C1(clknet_1_1__leaf_net859),
    .D1(net860),
    .X(net856));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net413),
    .A1(net289),
    .A2(net898),
    .A3(net850),
    .S0(clknet_1_0__leaf_net826),
    .S1(net365),
    .X(net414));
 sky130_fd_sc_hd__a2111o_1 c477 (.A1(net850),
    .A2(clknet_1_0__leaf_net403),
    .B1(net412),
    .C1(net693),
    .D1(net695),
    .X(net415));
 sky130_fd_sc_hd__a2111o_1 c478 (.A1(net409),
    .A2(net413),
    .B1(clknet_1_0__leaf_net386),
    .C1(net898),
    .D1(net694),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net288),
    .A1(net413),
    .A2(net291),
    .A3(clknet_1_1__leaf_net859),
    .S0(net679),
    .S1(net695),
    .X(net417));
 sky130_fd_sc_hd__sdfbbp_1 c480 (.CLK(clknet_2_3__leaf_clk),
    .D(net405),
    .RESET_B(net417),
    .SCD(net899),
    .SCE(clknet_1_0__leaf_net826),
    .SET_B(net694),
    .Q(net840));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net407),
    .A1(net416),
    .A2(net851),
    .A3(net169),
    .S0(net412),
    .S1(net694),
    .X(net418));
 sky130_fd_sc_hd__sdfbbn_1 c482 (.CLK_N(clknet_leaf_16_clk),
    .D(net885),
    .RESET_B(net415),
    .SCD(net412),
    .SCE(net692),
    .SET_B(net858),
    .Q(net420),
    .Q_N(net419));
 sky130_fd_sc_hd__and2_4 c504 (.A(net675),
    .B(net82),
    .X(net421));
 sky130_fd_sc_hd__and2_0 c505 (.A(net819),
    .B(net84),
    .X(net422));
 sky130_fd_sc_hd__and2_4 c506 (.A(net421),
    .B(net886),
    .X(net423));
 sky130_fd_sc_hd__and2_0 c507 (.A(net332),
    .B(net421),
    .X(net424));
 sky130_fd_sc_hd__and2_1 c508 (.A(net320),
    .B(net915),
    .X(net425));
 sky130_fd_sc_hd__and2_1 c509 (.A(net216),
    .B(net421),
    .X(net426));
 sky130_fd_sc_hd__and3_4 c510 (.A(net425),
    .B(net886),
    .C(net916),
    .X(net427));
 sky130_fd_sc_hd__sdfxtp_1 c511 (.CLK(clknet_leaf_32_clk),
    .D(net323),
    .SCD(net333),
    .SCE(net921),
    .Q(net428));
 sky130_fd_sc_hd__sdfxtp_4 c512 (.CLK(clknet_leaf_32_clk),
    .D(net921),
    .SCD(net319),
    .SCE(net425),
    .Q(net837));
 sky130_fd_sc_hd__dfbbn_1 c513 (.CLK_N(clknet_leaf_32_clk),
    .D(net426),
    .RESET_B(net886),
    .SET_B(net427),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__and2_2 c514 (.A(net425),
    .B(net423),
    .X(net431));
 sky130_fd_sc_hd__and2_1 c515 (.A(net424),
    .B(net837),
    .X(net432));
 sky130_fd_sc_hd__and3_1 c516 (.A(net431),
    .B(net202),
    .C(net886),
    .X(net433));
 sky130_fd_sc_hd__dfbbn_1 c517 (.CLK_N(clknet_leaf_32_clk),
    .D(net963),
    .RESET_B(net426),
    .SET_B(net318),
    .Q(net435),
    .Q_N(net434));
 sky130_fd_sc_hd__and2_4 c518 (.A(net206),
    .B(net424),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net435),
    .A1(net427),
    .A2(net436),
    .A3(net425),
    .S0(net431),
    .S1(net432),
    .X(net437));
 sky130_fd_sc_hd__mux4_2 c520 (.A0(net434),
    .A1(net317),
    .A2(net436),
    .A3(net837),
    .S0(net427),
    .S1(net886),
    .X(net438));
 sky130_fd_sc_hd__a2111o_1 c521 (.A1(net438),
    .A2(net431),
    .B1(net772),
    .C1(net887),
    .D1(net662),
    .X(net439));
 sky130_fd_sc_hd__mux4_2 c522 (.A0(net433),
    .A1(net437),
    .A2(net428),
    .A3(net427),
    .S0(net889),
    .S1(net886),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net427),
    .A1(net425),
    .A2(net880),
    .A3(net438),
    .S0(net436),
    .S1(net889),
    .X(net441));
 sky130_fd_sc_hd__dfbbp_1 c524 (.CLK(clknet_leaf_31_clk),
    .D(net441),
    .RESET_B(net438),
    .SET_B(net71),
    .Q(net442));
 sky130_fd_sc_hd__and3_1 c525 (.A(net342),
    .B(net431),
    .C(net886),
    .X(net443));
 sky130_fd_sc_hd__and2_4 c526 (.A(net912),
    .B(net832),
    .X(net444));
 sky130_fd_sc_hd__and2_0 c527 (.A(net431),
    .B(net355),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c528 (.A(net84),
    .B(net883),
    .C(net423),
    .X(net446));
 sky130_fd_sc_hd__dfstp_1 c529 (.CLK(clknet_leaf_32_clk),
    .D(net426),
    .SET_B(net446),
    .Q(net447));
 sky130_fd_sc_hd__and2_0 c530 (.A(net330),
    .B(net432),
    .X(net448));
 sky130_fd_sc_hd__and3_1 c531 (.A(net447),
    .B(net84),
    .C(net355),
    .X(net449));
 sky130_fd_sc_hd__and3_1 c532 (.A(net438),
    .B(net969),
    .C(net886),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c533 (.A0(net449),
    .A1(net233),
    .A2(net447),
    .A3(net348),
    .S0(net227),
    .S1(net444),
    .X(net451));
 sky130_fd_sc_hd__and3_4 c534 (.A(net338),
    .B(net69),
    .C(net423),
    .X(net452));
 sky130_fd_sc_hd__and2_0 c535 (.A(net886),
    .B(net339),
    .X(net453));
 sky130_fd_sc_hd__and2_0 c536 (.A(net450),
    .B(net313),
    .X(net454));
 sky130_fd_sc_hd__a2111o_4 c537 (.A1(net227),
    .A2(net825),
    .B1(net793),
    .C1(net880),
    .D1(net975),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net445),
    .A1(net452),
    .A2(net436),
    .A3(net444),
    .S0(net348),
    .S1(net770),
    .X(net456));
 sky130_fd_sc_hd__sdfstp_1 c539 (.CLK(clknet_leaf_32_clk),
    .D(net319),
    .SCD(net448),
    .SCE(net452),
    .SET_B(net926),
    .Q(net457));
 sky130_fd_sc_hd__sdfbbn_1 c540 (.CLK_N(clknet_leaf_36_clk),
    .D(net448),
    .RESET_B(net447),
    .SCD(net455),
    .SCE(net445),
    .SET_B(net319),
    .Q(net459),
    .Q_N(net458));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net453),
    .A1(net925),
    .A2(net438),
    .A3(net452),
    .S0(net444),
    .S1(net459),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net457),
    .A1(net779),
    .A2(net338),
    .A3(net313),
    .S0(net447),
    .S1(net348),
    .X(net461));
 sky130_fd_sc_hd__sdfbbp_1 c543 (.CLK(clknet_leaf_33_clk),
    .D(net461),
    .RESET_B(net455),
    .SCD(net432),
    .SCE(net431),
    .SET_B(net937),
    .Q(net463),
    .Q_N(net462));
 sky130_fd_sc_hd__sdfbbn_2 c544 (.CLK_N(clknet_leaf_33_clk),
    .D(net446),
    .RESET_B(net887),
    .SCD(net461),
    .SCE(net449),
    .SET_B(net699),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net214),
    .A1(net436),
    .A2(net453),
    .A3(net465),
    .S0(net792),
    .S1(net458),
    .X(net466));
 sky130_fd_sc_hd__dlrbn_1 c546 (.D(net83),
    .GATE_N(clknet_leaf_35_clk),
    .RESET_B(net444),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__dlrbn_1 c547 (.D(net311),
    .GATE_N(clknet_leaf_34_clk),
    .RESET_B(net969),
    .Q(net470),
    .Q_N(net469));
 sky130_fd_sc_hd__and2_0 c548 (.A(net469),
    .B(net945),
    .X(net471));
 sky130_fd_sc_hd__and3_2 c549 (.A(net355),
    .B(net459),
    .C(net436),
    .X(net472));
 sky130_fd_sc_hd__dlrbp_1 c550 (.D(clknet_1_1__leaf_net375),
    .GATE(clknet_leaf_35_clk),
    .RESET_B(net941),
    .Q(net473));
 sky130_fd_sc_hd__and2_2 c551 (.A(net800),
    .B(net355),
    .X(net474));
 sky130_fd_sc_hd__and3_2 c552 (.A(net471),
    .B(net450),
    .C(net458),
    .X(net475));
 sky130_fd_sc_hd__and3_2 c553 (.A(net459),
    .B(net470),
    .C(net800),
    .X(net476));
 sky130_fd_sc_hd__dlrbp_1 c554 (.D(net474),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(net911),
    .Q(net477));
 sky130_fd_sc_hd__and3_1 c555 (.A(net795),
    .B(net476),
    .C(net452),
    .X(net478));
 sky130_fd_sc_hd__sdfxbp_1 c556 (.CLK(clknet_leaf_35_clk),
    .D(clknet_1_1__leaf_net130),
    .SCD(net472),
    .SCE(net262),
    .Q(net479));
 sky130_fd_sc_hd__dlrtn_1 c557 (.D(net454),
    .GATE_N(clknet_leaf_34_clk),
    .RESET_B(net937),
    .Q(net480));
 sky130_fd_sc_hd__and3_2 c558 (.A(net477),
    .B(net480),
    .C(net377),
    .X(net829));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(net98),
    .A1(net263),
    .A2(net480),
    .A3(net825),
    .S0(net311),
    .S1(net472),
    .X(net481));
 sky130_fd_sc_hd__and3_1 c560 (.A(net478),
    .B(net480),
    .C(net701),
    .X(net482));
 sky130_fd_sc_hd__and2_0 c561 (.A(net482),
    .B(net701),
    .X(net483));
 sky130_fd_sc_hd__or4bb_2 c562 (.A(net473),
    .B(net467),
    .C_N(net880),
    .D_N(net701),
    .X(net484));
 sky130_fd_sc_hd__or4bb_2 c563 (.A(net470),
    .B(net476),
    .C_N(net837),
    .D_N(net701),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net480),
    .A1(net479),
    .A2(net482),
    .A3(net879),
    .S0(net484),
    .S1(net485),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net483),
    .A1(net450),
    .A2(net485),
    .A3(net98),
    .S0(net902),
    .S1(clknet_1_0__leaf_net702),
    .X(net487));
 sky130_fd_sc_hd__sdfbbn_1 c566 (.CLK_N(clknet_leaf_34_clk),
    .D(net263),
    .RESET_B(net487),
    .SCD(net443),
    .SCE(net476),
    .SET_B(clknet_1_1__leaf_net702),
    .Q(net488));
 sky130_fd_sc_hd__or4bb_1 c567 (.A(net391),
    .B(net377),
    .C_N(net465),
    .D_N(net988),
    .X(net489));
 sky130_fd_sc_hd__sedfxbp_1 c568 (.CLK(clknet_leaf_14_clk),
    .D(net484),
    .DE(net880),
    .SCD(net485),
    .SCE(clknet_1_0__leaf_net281),
    .Q(net490));
 sky130_fd_sc_hd__a2111o_1 c569 (.A1(net889),
    .A2(net485),
    .B1(net882),
    .C1(net150),
    .D1(net669),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net356),
    .A1(net472),
    .A2(net902),
    .A3(net391),
    .S0(net228),
    .S1(clknet_1_0__leaf_net281),
    .X(net492));
 sky130_fd_sc_hd__sdfbbp_1 c571 (.CLK(clknet_leaf_35_clk),
    .D(net489),
    .RESET_B(net356),
    .SCD(net895),
    .SCE(net467),
    .SET_B(net878),
    .Q(net494),
    .Q_N(net493));
 sky130_fd_sc_hd__sdfbbn_1 c572 (.CLK_N(clknet_leaf_34_clk),
    .D(net452),
    .RESET_B(net217),
    .SCD(clknet_1_0__leaf_net389),
    .SCE(net878),
    .SET_B(clknet_1_1__leaf_net655),
    .Q(net495));
 sky130_fd_sc_hd__a2111o_1 c573 (.A1(net468),
    .A2(net452),
    .B1(net889),
    .C1(net891),
    .D1(net356),
    .X(net496));
 sky130_fd_sc_hd__sdfbbn_1 c574 (.CLK_N(clknet_leaf_14_clk),
    .D(net485),
    .RESET_B(net12),
    .SCD(clknet_1_0__leaf_net281),
    .SCE(net377),
    .SET_B(net894),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net228),
    .A1(net825),
    .A2(net476),
    .A3(clknet_1_0__leaf_net389),
    .S0(net497),
    .S1(clknet_1_0__leaf_net386),
    .X(net499));
 sky130_fd_sc_hd__or4bb_4 c576 (.A(net151),
    .B(net356),
    .C_N(net829),
    .D_N(net465),
    .X(net500));
 sky130_fd_sc_hd__or4bb_4 c577 (.A(net399),
    .B(net488),
    .C_N(net468),
    .D_N(net496),
    .X(net501));
 sky130_fd_sc_hd__sdfbbp_1 c578 (.CLK(clknet_leaf_23_clk),
    .D(net446),
    .RESET_B(net385),
    .SCD(clknet_1_0__leaf_net501),
    .SCE(net900),
    .SET_B(net703),
    .Q(net503),
    .Q_N(net502));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net476),
    .A1(net496),
    .A2(net493),
    .A3(net502),
    .S0(clknet_1_0__leaf_net501),
    .S1(net894),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(clknet_1_0__leaf_net389),
    .A1(net446),
    .A2(net468),
    .A3(net503),
    .S0(net476),
    .S1(clknet_1_1__leaf_net655),
    .X(net505));
 sky130_fd_sc_hd__sdfbbn_1 c581 (.CLK_N(clknet_leaf_23_clk),
    .D(net950),
    .RESET_B(net377),
    .SCD(net837),
    .SCE(clknet_1_1__leaf_net501),
    .SET_B(net502),
    .Q(net506));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net506),
    .A1(net500),
    .A2(net377),
    .A3(clknet_1_1__leaf_net501),
    .S0(net502),
    .S1(clknet_1_0__leaf_net834),
    .X(net507));
 sky130_fd_sc_hd__sdfbbn_1 c583 (.CLK_N(clknet_leaf_23_clk),
    .D(net957),
    .RESET_B(net494),
    .SCD(net500),
    .SCE(net503),
    .SET_B(net475),
    .Q(net509),
    .Q_N(net508));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(clknet_1_0__leaf_net501),
    .A1(net505),
    .A2(net508),
    .A3(net890),
    .S0(net910),
    .S1(net476),
    .X(net510));
 sky130_fd_sc_hd__or4bb_1 c585 (.A(net503),
    .B(net476),
    .C_N(net704),
    .D_N(net705),
    .X(net511));
 sky130_fd_sc_hd__sdfbbp_1 c586 (.CLK(clknet_leaf_23_clk),
    .D(net371),
    .RESET_B(net511),
    .SCD(net825),
    .SCE(net502),
    .SET_B(clknet_1_1__leaf_net501),
    .Q(net512));
 sky130_fd_sc_hd__sdfbbn_1 c587 (.CLK_N(clknet_leaf_23_clk),
    .D(net960),
    .RESET_B(net503),
    .SCD(clknet_1_1__leaf_net501),
    .SCE(net511),
    .SET_B(net837),
    .Q(net513));
 sky130_fd_sc_hd__sdfbbn_1 c588 (.CLK_N(clknet_leaf_22_clk),
    .D(net224),
    .RESET_B(net24),
    .SCD(net462),
    .SCE(clknet_1_0__leaf_net826),
    .SET_B(net822),
    .Q(net515),
    .Q_N(net514));
 sky130_fd_sc_hd__sdfbbp_1 c589 (.CLK(clknet_leaf_14_clk),
    .D(net420),
    .RESET_B(net772),
    .SCD(net909),
    .SCE(net224),
    .SET_B(net829),
    .Q(net517),
    .Q_N(net516));
 sky130_fd_sc_hd__sdfbbn_1 c590 (.CLK_N(clknet_leaf_15_clk),
    .D(net472),
    .RESET_B(net517),
    .SCD(net829),
    .SCE(clknet_1_1__leaf_net299),
    .SET_B(net695),
    .Q(net518));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net12),
    .A1(clknet_1_0__leaf_net299),
    .A2(net902),
    .A3(clknet_1_0__leaf_net826),
    .S0(net779),
    .S1(net695),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net513),
    .A1(net516),
    .A2(net24),
    .A3(clknet_1_0__leaf_net826),
    .S0(net694),
    .S1(clknet_1_1__leaf_net834),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_0__leaf_net299),
    .A1(net464),
    .A2(net372),
    .A3(net691),
    .S0(net693),
    .S1(net694),
    .X(net521));
 sky130_fd_sc_hd__sdfbbn_1 c594 (.CLK_N(clknet_leaf_22_clk),
    .D(clknet_1_1__leaf_net299),
    .RESET_B(net372),
    .SCD(net514),
    .SCE(net24),
    .SET_B(net954),
    .Q(net523),
    .Q_N(net522));
 sky130_fd_sc_hd__sdfbbp_1 c595 (.CLK(clknet_leaf_15_clk),
    .D(net879),
    .RESET_B(net24),
    .SCD(clknet_1_1__leaf_net655),
    .SCE(net970),
    .SET_B(net708),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__a2111o_2 c596 (.A1(net524),
    .A2(net881),
    .B1(net706),
    .C1(net707),
    .D1(net708),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net463),
    .A1(net512),
    .A2(net829),
    .A3(clknet_1_1__leaf_net655),
    .S0(net695),
    .S1(net708),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net490),
    .A1(net420),
    .A2(net837),
    .A3(net464),
    .S0(net894),
    .S1(net695),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net518),
    .A1(net792),
    .A2(net825),
    .A3(net444),
    .S0(clknet_1_1__leaf_net655),
    .S1(net706),
    .X(net529));
 sky130_fd_sc_hd__a2111o_1 c600 (.A1(net527),
    .A2(net837),
    .B1(net694),
    .C1(net708),
    .D1(net709),
    .X(net530));
 sky130_fd_sc_hd__mux4_2 c601 (.A0(clknet_1_1__leaf_net403),
    .A1(net528),
    .A2(net837),
    .A3(net875),
    .S0(clknet_1_0__leaf_net834),
    .S1(net708),
    .X(net531));
 sky130_fd_sc_hd__sdfbbn_1 c602 (.CLK_N(clknet_leaf_16_clk),
    .D(clknet_1_1__leaf_net531),
    .RESET_B(net24),
    .SCD(net972),
    .SCE(net298),
    .SET_B(net962),
    .Q(net877),
    .Q_N(net532));
 sky130_fd_sc_hd__mux4_2 c603 (.A0(net882),
    .A1(net532),
    .A2(net875),
    .A3(net706),
    .S0(net707),
    .S1(net709),
    .X(net533));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_leaf_16_clk),
    .D(net772),
    .RESET_B(net902),
    .SCD(net986),
    .SCE(net533),
    .SET_B(net962),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net138),
    .A1(net533),
    .A2(clknet_1_0__leaf_net531),
    .A3(net532),
    .S0(net472),
    .S1(net692),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net530),
    .A1(net902),
    .A2(net534),
    .A3(net533),
    .S0(net709),
    .S1(net977),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net525),
    .A1(net877),
    .A2(net535),
    .A3(net779),
    .S0(net533),
    .S1(net977),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net534),
    .A1(net690),
    .A2(net695),
    .A3(net708),
    .S0(net710),
    .S1(net712),
    .X(net539));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net800),
    .A1(net798),
    .A2(net760),
    .A3(net818),
    .S0(net771),
    .S1(net802),
    .X(net0));
 sky130_fd_sc_hd__and2_0 c63 (.A(net798),
    .B(net895),
    .X(net1));
 sky130_fd_sc_hd__and2_0 c630 (.A(net71),
    .B(net886),
    .X(net540));
 sky130_fd_sc_hd__or4bb_1 c631 (.A(net428),
    .B(net770),
    .C_N(net436),
    .D_N(net922),
    .X(net541));
 sky130_fd_sc_hd__and2_1 c632 (.A(net541),
    .B(net884),
    .X(net542));
 sky130_fd_sc_hd__and2_0 c633 (.A(net541),
    .B(net542),
    .X(net543));
 sky130_fd_sc_hd__and2_0 c634 (.A(net202),
    .B(net917),
    .X(net544));
 sky130_fd_sc_hd__and2_1 c635 (.A(net430),
    .B(net69),
    .X(net545));
 sky130_fd_sc_hd__dlrtn_1 c636 (.D(net543),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net923),
    .Q(net546));
 sky130_fd_sc_hd__and2_1 c637 (.A(net544),
    .B(net542),
    .X(net547));
 sky130_fd_sc_hd__and2_2 c638 (.A(net544),
    .B(net918),
    .X(net548));
 sky130_fd_sc_hd__and3_1 c639 (.A(net442),
    .B(net540),
    .C(net887),
    .X(net549));
 sky130_fd_sc_hd__and2_1 c64 (.A(net813),
    .B(net4),
    .X(net2));
 sky130_fd_sc_hd__and2_2 c640 (.A(net318),
    .B(net542),
    .X(net550));
 sky130_fd_sc_hd__and2_1 c641 (.A(net548),
    .B(net542),
    .X(net551));
 sky130_fd_sc_hd__and2_1 c642 (.A(net542),
    .B(net919),
    .X(net552));
 sky130_fd_sc_hd__dlrtn_2 c643 (.D(net546),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net551),
    .Q(net553));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net549),
    .A1(net546),
    .A2(net553),
    .A3(net551),
    .S0(net548),
    .S1(net887),
    .X(net554));
 sky130_fd_sc_hd__and2_1 c645 (.A(net439),
    .B(net553),
    .X(net555));
 sky130_fd_sc_hd__sedfxbp_1 c646 (.CLK(clknet_leaf_29_clk),
    .D(net551),
    .DE(net880),
    .SCD(net553),
    .SCE(net966),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__or4bb_4 c647 (.A(net553),
    .B(net556),
    .C_N(net887),
    .D_N(net713),
    .X(net558));
 sky130_fd_sc_hd__or4bb_1 c648 (.A(net540),
    .B(net553),
    .C_N(net548),
    .D_N(net549),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net557),
    .A1(net559),
    .A2(net543),
    .A3(net551),
    .S0(net555),
    .S1(net558),
    .X(net560));
 sky130_fd_sc_hd__and2_4 c65 (.A(net820),
    .B(net903),
    .X(net3));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net437),
    .A1(net559),
    .A2(net551),
    .A3(net542),
    .S0(net69),
    .S1(net989),
    .X(net561));
 sky130_fd_sc_hd__or4bb_1 c651 (.A(net232),
    .B(net317),
    .C_N(net339),
    .D_N(net464),
    .X(net562));
 sky130_fd_sc_hd__and3_1 c652 (.A(net562),
    .B(net317),
    .C(net548),
    .X(net563));
 sky130_fd_sc_hd__or4bb_1 c653 (.A(net317),
    .B(net545),
    .C_N(net880),
    .D_N(net715),
    .X(net564));
 sky130_fd_sc_hd__sedfxtp_1 c654 (.CLK(clknet_leaf_30_clk),
    .D(net444),
    .DE(net887),
    .SCD(net563),
    .SCE(net981),
    .Q(net565));
 sky130_fd_sc_hd__and3_1 c655 (.A(net69),
    .B(net772),
    .C(net700),
    .X(net566));
 sky130_fd_sc_hd__sdfxbp_1 c656 (.CLK(clknet_leaf_29_clk),
    .D(net432),
    .SCD(net880),
    .SCE(net550),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__sedfxtp_2 c657 (.CLK(clknet_leaf_30_clk),
    .D(net564),
    .DE(net444),
    .SCD(net550),
    .SCE(net971),
    .Q(net569));
 sky130_fd_sc_hd__sedfxtp_4 c658 (.CLK(clknet_leaf_29_clk),
    .D(net563),
    .DE(net569),
    .SCD(net552),
    .SCE(net880),
    .Q(net570));
 sky130_fd_sc_hd__and3_2 c659 (.A(net569),
    .B(net570),
    .C(net567),
    .X(net571));
 sky130_fd_sc_hd__and2_4 c66 (.A(net810),
    .B(net895),
    .X(net4));
 sky130_fd_sc_hd__or4bb_1 c660 (.A(net339),
    .B(net566),
    .C_N(net571),
    .D_N(net697),
    .X(net572));
 sky130_fd_sc_hd__sdfrbp_1 c661 (.CLK(clknet_leaf_30_clk),
    .D(net958),
    .RESET_B(net555),
    .SCD(net548),
    .SCE(net339),
    .Q(net574),
    .Q_N(net573));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net552),
    .A1(net789),
    .A2(net568),
    .A3(net563),
    .S0(net571),
    .S1(net551),
    .X(net575));
 sky130_fd_sc_hd__a2111o_1 c663 (.A1(net423),
    .A2(net572),
    .B1(net570),
    .C1(net887),
    .D1(clknet_1_0__leaf_net716),
    .X(net576));
 sky130_fd_sc_hd__mux4_2 c664 (.A0(net574),
    .A1(net69),
    .A2(clknet_1_0__leaf_net576),
    .A3(net317),
    .S0(net571),
    .S1(net570),
    .X(net577));
 sky130_fd_sc_hd__sdfbbp_1 c665 (.CLK(clknet_leaf_30_clk),
    .D(net202),
    .RESET_B(clknet_1_0__leaf_net576),
    .SCD(net550),
    .SCE(net571),
    .SET_B(net573),
    .Q(net578));
 sky130_fd_sc_hd__or4bb_1 c666 (.A(net578),
    .B(net570),
    .C_N(net715),
    .D_N(clknet_1_0__leaf_net716),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(net348),
    .A1(net574),
    .A2(clknet_1_0__leaf_net577),
    .A3(net569),
    .S0(net563),
    .S1(clknet_1_0__leaf_net716),
    .X(net580));
 sky130_fd_sc_hd__sdfrbp_1 c668 (.CLK(clknet_leaf_29_clk),
    .D(net953),
    .RESET_B(net552),
    .SCD(net571),
    .SCE(net455),
    .Q(net581));
 sky130_fd_sc_hd__mux4_1 c669 (.A0(net579),
    .A1(net465),
    .A2(clknet_1_0__leaf_net580),
    .A3(net570),
    .S0(net569),
    .S1(net714),
    .X(net582));
 sky130_fd_sc_hd__and2_0 c67 (.A(net2),
    .B(net903),
    .X(net5));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(net227),
    .A1(net574),
    .A2(clknet_1_0__leaf_net580),
    .A3(net567),
    .S0(net920),
    .S1(net717),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net581),
    .A1(net571),
    .A2(net920),
    .A3(net573),
    .S0(clknet_1_0__leaf_net580),
    .S1(net718),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(net455),
    .A1(net547),
    .A2(clknet_1_0__leaf_net577),
    .A3(net931),
    .S0(net233),
    .S1(clknet_1_1__leaf_net580),
    .X(net585));
 sky130_fd_sc_hd__sdfrtn_1 c673 (.CLK_N(clknet_leaf_33_clk),
    .D(net547),
    .RESET_B(net558),
    .SCD(net772),
    .SCE(net890),
    .Q(net586));
 sky130_fd_sc_hd__or4bb_1 c674 (.A(net571),
    .B(net545),
    .C_N(net553),
    .D_N(net894),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net555),
    .A1(net474),
    .A2(net890),
    .A3(net233),
    .S0(net558),
    .S1(net653),
    .X(net588));
 sky130_fd_sc_hd__sdfrtp_4 c676 (.CLK(clknet_leaf_28_clk),
    .D(net558),
    .RESET_B(clknet_1_1__leaf_net580),
    .SCD(net890),
    .SCE(net721),
    .Q(net589));
 sky130_fd_sc_hd__buf_1 c677 (.A(net759),
    .X(net590));
 sky130_fd_sc_hd__buf_1 c678 (.A(net759),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(clknet_1_1__leaf_net580),
    .A1(net587),
    .A2(net890),
    .A3(net884),
    .S0(net880),
    .S1(net720),
    .X(net592));
 sky130_fd_sc_hd__or4bb_1 c68 (.A(net772),
    .B(net895),
    .C_N(net797),
    .D_N(net801),
    .X(net6));
 sky130_fd_sc_hd__and3_1 c680 (.A(net772),
    .B(net789),
    .C(net721),
    .X(net593));
 sky130_fd_sc_hd__and3_1 c681 (.A(net545),
    .B(net482),
    .C(net589),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(net558),
    .A1(net594),
    .A2(net793),
    .A3(net698),
    .S0(clknet_1_0__leaf_net716),
    .S1(net723),
    .X(net595));
 sky130_fd_sc_hd__sdfrtp_1 c683 (.CLK(clknet_leaf_24_clk),
    .D(net590),
    .RESET_B(net475),
    .SCD(net436),
    .SCE(net589),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net475),
    .A1(net596),
    .A2(net890),
    .A3(net548),
    .S0(net589),
    .S1(net723),
    .X(net597));
 sky130_fd_sc_hd__mux4_2 c685 (.A0(net436),
    .A1(net930),
    .A2(net590),
    .A3(net596),
    .S0(clknet_1_0__leaf_net577),
    .S1(net558),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net595),
    .A1(net596),
    .A2(net558),
    .A3(net589),
    .S0(net591),
    .S1(net719),
    .X(net599));
 sky130_fd_sc_hd__sdfxtp_1 c687 (.CLK(clknet_leaf_27_clk),
    .D(net599),
    .SCD(net973),
    .SCE(net725),
    .Q(net600));
 sky130_fd_sc_hd__or4bb_4 c688 (.A(net793),
    .B(net596),
    .C_N(net589),
    .D_N(net725),
    .X(net601));
 sky130_fd_sc_hd__mux4_2 c689 (.A0(net443),
    .A1(net594),
    .A2(net601),
    .A3(net593),
    .S0(net436),
    .S1(net722),
    .X(net602));
 sky130_fd_sc_hd__and3_4 c69 (.A(net5),
    .B(net895),
    .C(net2),
    .X(net7));
 sky130_fd_sc_hd__a2111o_1 c690 (.A1(net600),
    .A2(net594),
    .B1(net553),
    .C1(net700),
    .D1(net725),
    .X(net603));
 sky130_fd_sc_hd__a2111o_1 c691 (.A1(net553),
    .A2(net603),
    .B1(net590),
    .C1(net589),
    .D1(net601),
    .X(net604));
 sky130_fd_sc_hd__sdfbbn_1 c692 (.CLK_N(clknet_leaf_24_clk),
    .D(net604),
    .RESET_B(net591),
    .SCD(net233),
    .SCE(net601),
    .SET_B(net722),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net566),
    .A1(clknet_1_1__leaf_net576),
    .A2(net475),
    .A3(net902),
    .S0(net878),
    .S1(clknet_1_1__leaf_net281),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net878),
    .A1(net548),
    .A2(net474),
    .A3(net372),
    .S0(net879),
    .S1(net722),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net550),
    .A1(net566),
    .A2(clknet_1_1__leaf_net576),
    .A3(net884),
    .S0(net878),
    .S1(net727),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net593),
    .A1(net475),
    .A2(net500),
    .A3(net878),
    .S0(clknet_1_1__leaf_net577),
    .S1(net723),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net884),
    .A1(net902),
    .A2(net779),
    .A3(net590),
    .S0(net550),
    .S1(net723),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net590),
    .A1(net772),
    .A2(net770),
    .A3(clknet_1_1__leaf_net576),
    .S0(clknet_1_0__leaf_net716),
    .S1(net729),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_0__leaf_net576),
    .A1(net593),
    .A2(net500),
    .A3(clknet_1_0__leaf_net716),
    .S0(net726),
    .S1(net728),
    .X(net613));
 sky130_fd_sc_hd__and2_0 c70 (.A(net817),
    .B(net7),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net589),
    .A1(net890),
    .A2(net772),
    .A3(net878),
    .S0(clknet_1_1__leaf_net577),
    .S1(net474),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net3),
    .A1(net500),
    .A2(net878),
    .A3(net593),
    .S0(net566),
    .S1(net893),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net21),
    .A1(net589),
    .A2(net372),
    .A3(clknet_1_1__leaf_net577),
    .S0(net879),
    .S1(net730),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net281),
    .A1(net550),
    .A2(net601),
    .A3(net605),
    .S0(net724),
    .S1(net893),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net474),
    .A1(net613),
    .A2(clknet_1_0__leaf_net598),
    .A3(net593),
    .S0(net728),
    .S1(net731),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_1__leaf_net386),
    .A1(net879),
    .A2(clknet_1_1__leaf_net576),
    .A3(net893),
    .S0(net732),
    .S1(net734),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(clknet_1_1__leaf_net281),
    .A1(net233),
    .A2(net566),
    .A3(net727),
    .S0(net893),
    .S1(clknet_1_0__leaf_net735),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net279),
    .A1(net548),
    .A2(net890),
    .A3(net566),
    .S0(net900),
    .S1(net737),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net878),
    .A1(net444),
    .A2(net728),
    .A3(net893),
    .S0(net733),
    .S1(net738),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(clknet_1_1__leaf_net577),
    .A1(net500),
    .A2(net601),
    .A3(net878),
    .S0(clknet_1_1__leaf_net386),
    .S1(net731),
    .X(net623));
 sky130_fd_sc_hd__and2_2 c71 (.A(net4),
    .B(net895),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net491),
    .A1(net550),
    .A2(net815),
    .A3(net601),
    .S0(clknet_1_0__leaf_net736),
    .S1(net739),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net550),
    .A1(net602),
    .A2(net893),
    .A3(clknet_1_1__leaf_net735),
    .S0(net740),
    .S1(net741),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net612),
    .A1(net500),
    .A2(net731),
    .A3(net740),
    .S0(net741),
    .S1(net742),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net626),
    .A1(net884),
    .A2(net475),
    .A3(net733),
    .S0(net741),
    .S1(net742),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(clknet_1_0__leaf_net598),
    .A1(net523),
    .A2(net881),
    .A3(net879),
    .S0(net900),
    .S1(net743),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net880),
    .A1(net526),
    .A2(net883),
    .A3(net522),
    .S0(net743),
    .S1(net744),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net884),
    .A1(net233),
    .A2(net770),
    .A3(net779),
    .S0(clknet_1_1__leaf_net716),
    .S1(net893),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net465),
    .A1(net298),
    .A2(clknet_1_1__leaf_net386),
    .A3(net526),
    .S0(net884),
    .S1(net747),
    .X(net631));
 sky130_fd_sc_hd__mux4_2 c718 (.A0(net815),
    .A1(net9),
    .A2(clknet_1_1__leaf_net598),
    .A3(net884),
    .S0(clknet_1_0__leaf_net736),
    .S1(net746),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net386),
    .A1(net606),
    .A2(net523),
    .A3(net822),
    .S0(net602),
    .S1(net746),
    .X(net633));
 sky130_fd_sc_hd__or4bb_1 c72 (.A(net8),
    .B(net7),
    .C_N(net891),
    .D_N(net813),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net539),
    .A1(clknet_1_0__leaf_net632),
    .A2(net601),
    .A3(net9),
    .S0(clknet_1_1__leaf_net672),
    .S1(net746),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net444),
    .A1(clknet_1_0__leaf_net633),
    .A2(net233),
    .A3(clknet_1_1__leaf_net736),
    .S0(net743),
    .S1(net744),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net298),
    .A1(net535),
    .A2(net515),
    .A3(net601),
    .S0(clknet_1_1__leaf_net386),
    .S1(net744),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net601),
    .A1(net602),
    .A2(net372),
    .A3(net822),
    .S0(net539),
    .S1(clknet_1_1__leaf_net716),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net535),
    .A1(net464),
    .A2(net653),
    .A3(clknet_1_1__leaf_net716),
    .S0(net743),
    .S1(net746),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net372),
    .A1(net634),
    .A2(net770),
    .A3(net9),
    .S0(net747),
    .S1(net749),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net526),
    .A1(net602),
    .A2(net70),
    .A3(net233),
    .S0(net745),
    .S1(net747),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net602),
    .A1(net881),
    .A2(net526),
    .A3(net893),
    .S0(net746),
    .S1(net967),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net515),
    .A1(clknet_1_1__leaf_net632),
    .A2(net822),
    .A3(net526),
    .S0(net743),
    .S1(net748),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net637),
    .A1(net881),
    .A2(net605),
    .A3(clknet_1_1__leaf_net672),
    .S0(net893),
    .S1(net743),
    .X(net643));
 sky130_fd_sc_hd__and2_1 c73 (.A(net8),
    .B(net801),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net879),
    .A1(net606),
    .A2(net514),
    .A3(clknet_1_1__leaf_net633),
    .S0(net711),
    .S1(net751),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net606),
    .A1(clknet_1_0__leaf_net633),
    .A2(clknet_1_1__leaf_net716),
    .A3(net893),
    .S0(net746),
    .S1(net749),
    .X(net645));
 sky130_fd_sc_hd__mux4_2 c732 (.A0(clknet_1_1__leaf_net386),
    .A1(clknet_1_0__leaf_net632),
    .A2(net747),
    .A3(net752),
    .S0(net754),
    .S1(net755),
    .X(net646));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(clknet_1_1__leaf_net646),
    .A1(net879),
    .A2(net881),
    .A3(net747),
    .S0(net756),
    .S1(net757),
    .X(net647));
 sky130_fd_sc_hd__mux4_2 c734 (.A0(clknet_1_1__leaf_net633),
    .A1(net638),
    .A2(clknet_1_0__leaf_net646),
    .A3(net747),
    .S0(net753),
    .S1(net758),
    .X(net648));
 sky130_fd_sc_hd__and2_2 c74 (.A(net891),
    .B(net7),
    .X(net12));
 sky130_fd_sc_hd__and3_4 c75 (.A(net10),
    .B(net891),
    .C(net895),
    .X(net13));
 sky130_fd_sc_hd__and2_0 c76 (.A(net12),
    .B(net891),
    .X(net14));
 sky130_fd_sc_hd__and2_0 c77 (.A(net10),
    .B(net13),
    .X(net15));
 sky130_fd_sc_hd__a2111o_4 c78 (.A1(net13),
    .A2(net15),
    .B1(net5),
    .C1(net895),
    .D1(net820),
    .X(net16));
 sky130_fd_sc_hd__and2_1 c79 (.A(net13),
    .B(net11),
    .X(net17));
 sky130_fd_sc_hd__a2111o_1 c80 (.A1(net16),
    .A2(net818),
    .B1(net15),
    .C1(net798),
    .D1(net12),
    .X(net18));
 sky130_fd_sc_hd__a2111o_2 c81 (.A1(net806),
    .A2(net7),
    .B1(net762),
    .C1(net14),
    .D1(net4),
    .X(net19));
 sky130_fd_sc_hd__and2_0 c82 (.A(net19),
    .B(net17),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c83 (.A0(net14),
    .A1(net7),
    .A2(net20),
    .A3(net19),
    .S0(net16),
    .S1(net13),
    .X(net21));
 sky130_fd_sc_hd__and2_2 c84 (.A(net801),
    .B(net2),
    .X(net22));
 sky130_fd_sc_hd__and3_1 c85 (.A(net19),
    .B(net761),
    .C(net16),
    .X(net23));
 sky130_fd_sc_hd__and2_4 c86 (.A(net16),
    .B(net22),
    .X(net24));
 sky130_fd_sc_hd__or4bb_4 c87 (.A(net24),
    .B(net2),
    .C_N(net22),
    .D_N(net19),
    .X(net25));
 sky130_fd_sc_hd__and2_0 c88 (.A(net814),
    .B(net11),
    .X(net26));
 sky130_fd_sc_hd__and3_2 c89 (.A(net26),
    .B(net797),
    .C(net24),
    .X(net27));
 sky130_fd_sc_hd__and2_4 c90 (.A(net25),
    .B(net23),
    .X(net28));
 sky130_fd_sc_hd__or4bb_1 c91 (.A(net2),
    .B(net23),
    .C_N(net28),
    .D_N(net4),
    .X(net29));
 sky130_fd_sc_hd__and2_1 c92 (.A(net762),
    .B(net22),
    .X(net30));
 sky130_fd_sc_hd__and2_2 c93 (.A(net25),
    .B(net24),
    .X(net31));
 sky130_fd_sc_hd__or4bb_1 c94 (.A(net30),
    .B(net4),
    .C_N(net24),
    .D_N(net797),
    .X(net32));
 sky130_fd_sc_hd__or4bb_1 c95 (.A(net32),
    .B(net992),
    .C_N(net23),
    .D_N(net26),
    .X(net33));
 sky130_fd_sc_hd__or4bb_1 c96 (.A(net32),
    .B(net31),
    .C_N(net27),
    .D_N(net992),
    .X(net34));
 sky130_fd_sc_hd__or4bb_1 c97 (.A(net26),
    .B(net19),
    .C_N(net803),
    .D_N(net11),
    .X(net35));
 sky130_fd_sc_hd__and2_1 c98 (.A(net23),
    .B(net28),
    .X(net36));
 sky130_fd_sc_hd__and3_1 c99 (.A(net33),
    .B(net32),
    .C(net31),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 merge740 (.A0(net570),
    .A1(net589),
    .A2(net547),
    .A3(net586),
    .S0(net474),
    .S1(net699),
    .X(net649));
 sky130_fd_sc_hd__dfxbp_1 s741 (.CLK(clknet_leaf_7_clk),
    .D(net39),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dfxbp_2 s742 (.CLK(clknet_leaf_7_clk),
    .D(net41),
    .Q(net867),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxtp_1 s743 (.CLK(clknet_leaf_8_clk),
    .D(net65),
    .Q(net854));
 sky130_fd_sc_hd__dfxtp_1 s744 (.CLK(clknet_leaf_8_clk),
    .D(net66),
    .Q(net847));
 sky130_fd_sc_hd__dfxtp_2 s745 (.CLK(clknet_leaf_43_clk),
    .D(net126),
    .Q(net653));
 sky130_fd_sc_hd__dlclkp_1 s746 (.CLK(clknet_leaf_43_clk),
    .GATE(net129),
    .GCLK(net859));
 sky130_fd_sc_hd__dlclkp_2 s747 (.CLK(clknet_leaf_43_clk),
    .GATE(net146),
    .GCLK(net654));
 sky130_fd_sc_hd__dlclkp_4 s748 (.CLK(clknet_leaf_4_clk),
    .GATE(net152),
    .GCLK(net655));
 sky130_fd_sc_hd__dlxbn_1 s749 (.D(net153),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net657),
    .Q_N(net656));
 sky130_fd_sc_hd__dlxbn_1 s750 (.D(net177),
    .GATE_N(clknet_leaf_6_clk),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dlxbp_1 s751 (.D(net178),
    .GATE(clknet_leaf_10_clk),
    .Q(net869),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxtn_2 s752 (.D(net179),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net875));
 sky130_fd_sc_hd__dlxtn_1 s753 (.D(net189),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net661));
 sky130_fd_sc_hd__dlxtn_1 s754 (.D(net197),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net828));
 sky130_fd_sc_hd__dlxtp_1 s755 (.D(net218),
    .GATE(clknet_leaf_40_clk),
    .Q(net662));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s756 (.D(net261),
    .SLEEP_B(clknet_leaf_0_clk),
    .Q(net663));
 sky130_fd_sc_hd__dfxbp_1 s757 (.CLK(clknet_leaf_1_clk),
    .D(net269),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfxbp_1 s758 (.CLK(clknet_leaf_3_clk),
    .D(net278),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfxtp_1 s759 (.CLK(clknet_leaf_3_clk),
    .D(net284),
    .Q(net668));
 sky130_fd_sc_hd__dfxtp_1 s760 (.CLK(clknet_leaf_2_clk),
    .D(net285),
    .Q(net669));
 sky130_fd_sc_hd__dfxtp_1 s761 (.CLK(clknet_leaf_3_clk),
    .D(net294),
    .Q(net670));
 sky130_fd_sc_hd__dlclkp_1 s762 (.CLK(clknet_leaf_12_clk),
    .GATE(net302),
    .GCLK(net671));
 sky130_fd_sc_hd__dlclkp_2 s763 (.CLK(clknet_leaf_13_clk),
    .GATE(net305),
    .GCLK(net672));
 sky130_fd_sc_hd__dlclkp_4 s764 (.CLK(clknet_leaf_11_clk),
    .GATE(net306),
    .GCLK(net868));
 sky130_fd_sc_hd__dlxbn_1 s765 (.D(net307),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net870),
    .Q_N(net865));
 sky130_fd_sc_hd__dlxbn_1 s766 (.D(net308),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net866),
    .Q_N(net673));
 sky130_fd_sc_hd__dlxbp_1 s767 (.D(net309),
    .GATE(clknet_leaf_10_clk),
    .Q(net864),
    .Q_N(net674));
 sky130_fd_sc_hd__dlxtn_2 s768 (.D(net329),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net675));
 sky130_fd_sc_hd__dlxtn_1 s769 (.D(net331),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net676));
 sky130_fd_sc_hd__dlxtn_1 s770 (.D(net334),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net677));
 sky130_fd_sc_hd__dlxtp_1 s771 (.D(net341),
    .GATE(clknet_leaf_37_clk),
    .Q(net678));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s772 (.D(net343),
    .SLEEP_B(clknet_leaf_36_clk),
    .Q(net679));
 sky130_fd_sc_hd__dfxbp_1 s773 (.CLK(clknet_leaf_36_clk),
    .D(net357),
    .Q(net680));
 sky130_fd_sc_hd__dfxbp_1 s774 (.CLK(clknet_leaf_1_clk),
    .D(net362),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dfxtp_1 s775 (.CLK(clknet_leaf_36_clk),
    .D(net374),
    .Q(net683));
 sky130_fd_sc_hd__dfxtp_1 s776 (.CLK(clknet_leaf_35_clk),
    .D(net376),
    .Q(net684));
 sky130_fd_sc_hd__dfxtp_1 s777 (.CLK(clknet_leaf_35_clk),
    .D(net378),
    .Q(net685));
 sky130_fd_sc_hd__dlclkp_1 s778 (.CLK(clknet_leaf_35_clk),
    .GATE(net379),
    .GCLK(net686));
 sky130_fd_sc_hd__dlclkp_2 s779 (.CLK(clknet_leaf_2_clk),
    .GATE(net384),
    .GCLK(net687));
 sky130_fd_sc_hd__dlclkp_4 s780 (.CLK(clknet_leaf_14_clk),
    .GATE(net392),
    .GCLK(net688));
 sky130_fd_sc_hd__dlxbn_1 s781 (.D(net394),
    .GATE_N(clknet_leaf_14_clk),
    .Q(net689));
 sky130_fd_sc_hd__dlxbn_1 s782 (.D(net398),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net691),
    .Q_N(net690));
 sky130_fd_sc_hd__dlxbp_1 s783 (.D(net402),
    .GATE(clknet_leaf_15_clk),
    .Q(net693),
    .Q_N(net692));
 sky130_fd_sc_hd__dlxtn_2 s784 (.D(net406),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net694));
 sky130_fd_sc_hd__dlxtn_1 s785 (.D(net410),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net848));
 sky130_fd_sc_hd__dlxtn_1 s786 (.D(net411),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net860));
 sky130_fd_sc_hd__dlxtp_1 s787 (.D(net414),
    .GATE(clknet_leaf_14_clk),
    .Q(net695));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s788 (.D(net418),
    .SLEEP_B(clknet_leaf_16_clk),
    .Q(net858));
 sky130_fd_sc_hd__dfxbp_1 s789 (.CLK(clknet_leaf_33_clk),
    .D(net451),
    .Q(net696));
 sky130_fd_sc_hd__dfxbp_1 s790 (.CLK(clknet_leaf_33_clk),
    .D(net456),
    .Q(net698),
    .Q_N(net697));
 sky130_fd_sc_hd__dfxtp_1 s791 (.CLK(clknet_leaf_33_clk),
    .D(net460),
    .Q(net699));
 sky130_fd_sc_hd__dfxtp_1 s792 (.CLK(clknet_leaf_33_clk),
    .D(net466),
    .Q(net700));
 sky130_fd_sc_hd__dfxtp_1 s793 (.CLK(clknet_leaf_34_clk),
    .D(net481),
    .Q(net701));
 sky130_fd_sc_hd__dlclkp_1 s794 (.CLK(clknet_leaf_34_clk),
    .GATE(net486),
    .GCLK(net702));
 sky130_fd_sc_hd__dlclkp_2 s795 (.CLK(clknet_leaf_23_clk),
    .GATE(net492),
    .GCLK(net834));
 sky130_fd_sc_hd__dlclkp_4 s796 (.CLK(clknet_leaf_23_clk),
    .GATE(net499),
    .GCLK(net703));
 sky130_fd_sc_hd__dlxbn_1 s797 (.D(net504),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net704));
 sky130_fd_sc_hd__dlxbn_1 s798 (.D(net507),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net705));
 sky130_fd_sc_hd__dlxbp_1 s799 (.D(net510),
    .GATE(clknet_leaf_26_clk),
    .Q(net824));
 sky130_fd_sc_hd__dlxtn_1 s800 (.D(net519),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net706));
 sky130_fd_sc_hd__dlxtn_1 s801 (.D(net520),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net707));
 sky130_fd_sc_hd__dlxtn_2 s802 (.D(net521),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net708));
 sky130_fd_sc_hd__dlxtp_1 s803 (.D(net529),
    .GATE(clknet_leaf_15_clk),
    .Q(net709));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s804 (.D(net536),
    .SLEEP_B(clknet_leaf_16_clk),
    .Q(net710));
 sky130_fd_sc_hd__dfxbp_1 s805 (.CLK(clknet_leaf_18_clk),
    .D(net537),
    .Q(net711));
 sky130_fd_sc_hd__dfxbp_1 s806 (.CLK(clknet_leaf_18_clk),
    .D(net538),
    .Q(net712));
 sky130_fd_sc_hd__dfxtp_1 s807 (.CLK(clknet_leaf_31_clk),
    .D(net554),
    .Q(net713));
 sky130_fd_sc_hd__dfxtp_1 s808 (.CLK(clknet_leaf_30_clk),
    .D(net560),
    .Q(net714));
 sky130_fd_sc_hd__dfxtp_1 s809 (.CLK(clknet_leaf_30_clk),
    .D(net561),
    .Q(net715));
 sky130_fd_sc_hd__dlclkp_1 s810 (.CLK(clknet_leaf_29_clk),
    .GATE(net575),
    .GCLK(net716));
 sky130_fd_sc_hd__dlclkp_2 s811 (.CLK(clknet_leaf_29_clk),
    .GATE(net582),
    .GCLK(net717));
 sky130_fd_sc_hd__dlclkp_4 s812 (.CLK(clknet_leaf_28_clk),
    .GATE(net583),
    .GCLK(net718));
 sky130_fd_sc_hd__dlxbn_1 s813 (.D(net584),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net719));
 sky130_fd_sc_hd__dlxbn_1 s814 (.D(net585),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlxbp_1 s815 (.D(net588),
    .GATE(clknet_leaf_24_clk),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dlxtn_1 s816 (.D(net592),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net724));
 sky130_fd_sc_hd__dlxtn_1 s817 (.D(net597),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net725));
 sky130_fd_sc_hd__dlxtn_1 s818 (.D(net607),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net726));
 sky130_fd_sc_hd__dlxtp_1 s819 (.D(net608),
    .GATE(clknet_leaf_24_clk),
    .Q(net727));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s820 (.D(net609),
    .SLEEP_B(clknet_leaf_24_clk),
    .Q(net728));
 sky130_fd_sc_hd__dfxbp_1 s821 (.CLK(clknet_leaf_26_clk),
    .D(net610),
    .Q(net729));
 sky130_fd_sc_hd__dfxbp_1 s822 (.CLK(clknet_leaf_27_clk),
    .D(net611),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_1 s823 (.CLK(clknet_leaf_26_clk),
    .D(net614),
    .Q(net731));
 sky130_fd_sc_hd__dfxtp_1 s824 (.CLK(clknet_leaf_21_clk),
    .D(net615),
    .Q(net732));
 sky130_fd_sc_hd__dfxtp_1 s825 (.CLK(clknet_leaf_26_clk),
    .D(net616),
    .Q(net733));
 sky130_fd_sc_hd__dlclkp_1 s826 (.CLK(clknet_leaf_25_clk),
    .GATE(net617),
    .GCLK(net734));
 sky130_fd_sc_hd__dlclkp_2 s827 (.CLK(clknet_leaf_25_clk),
    .GATE(net618),
    .GCLK(net735));
 sky130_fd_sc_hd__dlclkp_4 s828 (.CLK(clknet_leaf_20_clk),
    .GATE(net619),
    .GCLK(net736));
 sky130_fd_sc_hd__dlxbn_1 s829 (.D(net620),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net737));
 sky130_fd_sc_hd__dlxbn_1 s830 (.D(net621),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net738));
 sky130_fd_sc_hd__dlxbp_1 s831 (.D(net622),
    .GATE(clknet_leaf_25_clk),
    .Q(net739));
 sky130_fd_sc_hd__dlxtn_1 s832 (.D(net623),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net740));
 sky130_fd_sc_hd__dlxtn_1 s833 (.D(net624),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s834 (.D(net625),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtp_1 s835 (.D(net627),
    .GATE(clknet_leaf_20_clk),
    .Q(net743));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s836 (.D(net628),
    .SLEEP_B(clknet_leaf_21_clk),
    .Q(net744));
 sky130_fd_sc_hd__dfxbp_1 s837 (.CLK(clknet_leaf_22_clk),
    .D(net629),
    .Q(net745));
 sky130_fd_sc_hd__dfxbp_2 s838 (.CLK(clknet_leaf_19_clk),
    .D(net630),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dfxtp_1 s839 (.CLK(clknet_leaf_18_clk),
    .D(net631),
    .Q(net748));
 sky130_fd_sc_hd__dfxtp_1 s840 (.CLK(clknet_leaf_19_clk),
    .D(net635),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_1 s841 (.CLK(clknet_leaf_22_clk),
    .D(net636),
    .Q(net750));
 sky130_fd_sc_hd__dlclkp_1 s842 (.CLK(clknet_leaf_19_clk),
    .GATE(net639),
    .GCLK(net751));
 sky130_fd_sc_hd__dlclkp_2 s843 (.CLK(clknet_leaf_18_clk),
    .GATE(net640),
    .GCLK(net752));
 sky130_fd_sc_hd__dlclkp_4 s844 (.CLK(clknet_leaf_19_clk),
    .GATE(net641),
    .GCLK(net753));
 sky130_fd_sc_hd__dlxbn_1 s845 (.D(net642),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net754));
 sky130_fd_sc_hd__dlxbn_1 s846 (.D(net643),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net823));
 sky130_fd_sc_hd__dlxbp_1 s847 (.D(net644),
    .GATE(clknet_leaf_19_clk),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dlxtn_1 s848 (.D(net645),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net757));
 sky130_fd_sc_hd__dlxtn_1 s849 (.D(net647),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net758));
 sky130_fd_sc_hd__dlxtn_4 s850 (.D(net648),
    .GATE_N(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dlxtp_1 s851 (.D(net649),
    .GATE(clknet_leaf_28_clk),
    .Q(net759));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(in0),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net761));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net762));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net763));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input6 (.A(in13),
    .X(net765));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in15),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net769));
 sky130_fd_sc_hd__buf_4 input11 (.A(in18),
    .X(net770));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net771));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net773));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net774));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_8 input20 (.A(in26),
    .X(net779));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(in27),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in28),
    .X(net781));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in3),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net784));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(in31),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net786));
 sky130_fd_sc_hd__buf_2 input28 (.A(in33),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net788));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net789));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net790));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net791));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net792));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net793));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net794));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net797));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net800));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net801));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(in5),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in50),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net807));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(in54),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in55),
    .X(net811));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(in57),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in58),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(in6),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net817));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net818));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net819));
 sky130_fd_sc_hd__buf_2 input61 (.A(in8),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in9),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net822),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net823),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net824),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net825),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(clknet_1_1__leaf_net826),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net827),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net828),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net829),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net830),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(clknet_1_1__leaf_net831),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net832),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net833),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(clknet_1_1__leaf_net834),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net835),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net836),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output78 (.A(net837),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net838),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output80 (.A(net839),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net840),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net841),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output83 (.A(net842),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net843),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net844),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net899),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net846),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net847),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net848),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net849),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net850),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net851),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net852),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net853),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net854),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net855),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net856),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net857),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net858),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(clknet_1_1__leaf_net859),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net860),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net861),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net862),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net863),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net864),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net865),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net866),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net867),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net868),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net869),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net870),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(clknet_1_1__leaf_net871),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net872),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output114 (.A(net873),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_1__leaf_net874),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net875),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output117 (.A(net876),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net877),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net491),
    .X(net878));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net842),
    .X(net879));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net904),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net440),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net138),
    .X(net882));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(net211),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net211),
    .X(net884));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net102),
    .X(net885));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(net422),
    .X(net887));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net199),
    .X(net888));
 sky130_fd_sc_hd__buf_4 fanout130 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net314),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net9),
    .X(net891));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net140),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net731),
    .X(net893));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net653),
    .X(net894));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net3),
    .X(net895));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net898),
    .X(net896));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout138 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net845),
    .X(net899));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(net70),
    .X(net900));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net857),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net815),
    .X(net902));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(net807),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net646 (.A(net646),
    .X(clknet_0_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_0__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net646 (.A(clknet_0_net646),
    .X(clknet_1_1__leaf_net646));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net736 (.A(net736),
    .X(clknet_0_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_0__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_1__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net632 (.A(net632),
    .X(clknet_0_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_0__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net632 (.A(clknet_0_net632),
    .X(clknet_1_1__leaf_net632));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net735 (.A(net735),
    .X(clknet_0_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_0__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net735 (.A(clknet_0_net735),
    .X(clknet_1_1__leaf_net735));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net716 (.A(net716),
    .X(clknet_0_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net716 (.A(clknet_0_net716),
    .X(clknet_1_1__leaf_net716));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net576 (.A(net576),
    .X(clknet_0_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net576 (.A(clknet_0_net576),
    .X(clknet_1_0__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net576 (.A(net924),
    .X(clknet_1_1__leaf_net576));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net598 (.A(net598),
    .X(clknet_0_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_0__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_1__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net834 (.A(net834),
    .X(clknet_0_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_0__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net834 (.A(clknet_0_net834),
    .X(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net531 (.A(net531),
    .X(clknet_0_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_0__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_1__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net826 (.A(net826),
    .X(clknet_0_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net826 (.A(clknet_0_net826),
    .X(clknet_1_1__leaf_net826));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net687 (.A(net687),
    .X(clknet_0_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_0__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net687 (.A(clknet_0_net687),
    .X(clknet_1_1__leaf_net687));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net846 (.A(net846),
    .X(clknet_0_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_1__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net386 (.A(net386),
    .X(clknet_0_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net386 (.A(clknet_0_net386),
    .X(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net633 (.A(net633),
    .X(clknet_0_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_0__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net633 (.A(clknet_0_net633),
    .X(clknet_1_1__leaf_net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net393 (.A(net393),
    .X(clknet_0_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_0__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net393 (.A(clknet_0_net393),
    .X(clknet_1_1__leaf_net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net686 (.A(net686),
    .X(clknet_0_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_0__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_1__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net672 (.A(net672),
    .X(clknet_0_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_0__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net672 (.A(clknet_0_net672),
    .X(clknet_1_1__leaf_net672));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net403 (.A(net403),
    .X(clknet_0_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_0__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net403 (.A(clknet_0_net403),
    .X(clknet_1_1__leaf_net403));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net831 (.A(net831),
    .X(clknet_0_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net831 (.A(clknet_0_net831),
    .X(clknet_1_0__leaf_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net831 (.A(clknet_0_net831),
    .X(clknet_1_1__leaf_net831));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net871 (.A(net871),
    .X(clknet_0_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_0__leaf_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net871 (.A(clknet_0_net871),
    .X(clknet_1_1__leaf_net871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net671 (.A(net671),
    .X(clknet_0_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_0__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net671 (.A(clknet_0_net671),
    .X(clknet_1_1__leaf_net671));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net154 (.A(net154),
    .X(clknet_0_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_0__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_1__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net855 (.A(net855),
    .X(clknet_0_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_0__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net855 (.A(clknet_0_net855),
    .X(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net859 (.A(net859),
    .X(clknet_0_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net874 (.A(net874),
    .X(clknet_0_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_0__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_1__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net155 (.A(net155),
    .X(clknet_0_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_0__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net155 (.A(clknet_0_net155),
    .X(clknet_1_1__leaf_net155));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net375 (.A(net375),
    .X(clknet_0_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_0__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net375 (.A(clknet_0_net375),
    .X(clknet_1_1__leaf_net375));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer1 (.A(net440),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net102),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net905),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net217),
    .X(net907));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer5 (.A(net907),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net217),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net217),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net910),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net85),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net28),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net913),
    .X(net914));
 sky130_fd_sc_hd__buf_2 rebuffer12 (.A(net675),
    .X(net915));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer13 (.A(net915),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net916),
    .X(net917));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer15 (.A(net917),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net918),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net423),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net423),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net423),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net922),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(clknet_0_net576),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net450),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net925),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net92),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer25 (.A(net927),
    .X(net928));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer26 (.A(net928),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net482),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net930),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net215),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net678),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net803),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net339),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net260),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net699),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net679),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net55),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net42),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net469),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net323),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net322),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net124),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net685),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net123),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net171),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net349),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net166),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net498),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net325),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net344),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net568),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net707),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net363),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net303),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net495),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net565),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net400),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net509),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net324),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net708),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net429),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net321),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net192),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net713),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net750),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net297),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net447),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net693),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net715),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net419),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net596),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net387),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net696),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net143),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net710),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net854),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net684),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net651),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net714),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net340),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net667),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net650),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net255),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net877),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net316),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net669),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net714),
    .X(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_RESET_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_D (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_D_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Q_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Q (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C_N (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_SCE (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_D1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_RESET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SET_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_Q (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_Q (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_SCE (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_SCD (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SCE (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_D_N (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_C (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_C (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_SCE (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Q (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_RESET_B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_C_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCE (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_SCD (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Q (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_SCE (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_S0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_RESET_B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCD (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A3 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_S0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCE (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SET_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Q (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_SCE (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Q (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_C_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_C (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_RESET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_RESET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_RESET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCD (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_SCD (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_SET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_C_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_RESET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_X (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_C_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_SCE (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_SCE (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_C1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A3 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_SET_B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCE (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_SCD (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCE (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A3 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_D_N (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_SET_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_RESET_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_X (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_S0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_Q (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SET_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_SET_B (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCD (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_C_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_Q (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_S1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_RESET_B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A0 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_D (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_RESET_B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_RESET_B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_D (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_Q (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_D (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_RESET_B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_RESET_B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SCE (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_D (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_C (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_C (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_B (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_X (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_SCD (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_C_N (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_C (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_X (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_DE (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_D (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_RESET_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_S1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_X (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_SET_B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_SCE (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_RESET_B (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCD (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_X (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCD (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q_N (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_Q (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_D_N (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Q_N (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_D_N (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_C_N (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Q (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_D (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_S1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge740_S0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_RESET_B (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SET_B (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_X (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_SCE (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCD (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SCD (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_SCD (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_C (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_C_N (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_X (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_SCD (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_SCD (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_SCE (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_X (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_B1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_C_N (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_SCD (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_Q (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_D (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_RESET_B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_X (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_D1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_X (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_S1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s745_Q (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_s772_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_C1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_S0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_C (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_s787_Q (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SET_B (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_D1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_SET_B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_Q (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_D1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_D1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_RESET_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_RESET_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_RESET_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_D_N (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_C_N (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_C (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_C (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_C (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_SCD (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_RESET_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_B1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_D1 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A0 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_C1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_SCE (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_C_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_D_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_D1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCE (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_D_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_C (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_D1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_SCE (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_D_N (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_C_N (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_C (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C_N (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_SCE (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SCE (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_D1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_C_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_D1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SET_B (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SCD (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_SET_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_SET_B (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_SCD (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SET_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C_N (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_RESET_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_SET_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_SET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_SCD (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_C_N (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_Q (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net859_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_s746_GCLK (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_s742_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_s752_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_D1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_SCE (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCD (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_DE (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C_N (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_C1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_SCE (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_SCD (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_C_N (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_DE (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_B1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S0 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_C (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_C1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_D1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_S1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_C (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_D (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_SET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_RESET_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_C1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_DE (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_C_N (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_C (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_C1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCE (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_D1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_SCE (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_SET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_SET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_B1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_SCE (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SCE (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_SET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_SCE (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_SCD (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_C_N (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_SCE (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_C1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_SCD (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_SCD (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_SET_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_D_N (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_D1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SCD (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_C1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_C (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C_N (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCD (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_SCE (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_C (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_SCE (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_C (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_C_N (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_D1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_SCD (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_D (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SCE (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_S0 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_RESET_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_D1 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_D_N (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net716_X (.DIODE(clknet_1_0__leaf_net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net834_X (.DIODE(clknet_1_1__leaf_net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_SCE (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCE (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net826_X (.DIODE(clknet_1_0__leaf_net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_D_N (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_RESET_B (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_C (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net386_X (.DIODE(clknet_1_0__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B1 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net386_X (.DIODE(clknet_1_1__leaf_net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S0 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net655_X (.DIODE(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_SET_B (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_SCD (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net655_X (.DIODE(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net855_X (.DIODE(clknet_1_1__leaf_net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_C (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_SET_B (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net859_X (.DIODE(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_D_N (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_C1 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net859_X (.DIODE(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_D_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_C (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SCD (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCE (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net792));
 sky130_fd_sc_hd__and2_1 clone1 (.A(net992),
    .B(net22),
    .X(net990));
 sky130_fd_sc_hd__and2_1 clone2 (.A(net82),
    .B(net81),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net16),
    .X(net992));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
