module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net617;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net664;
 wire clknet_1_0__leaf_net664;
 wire clknet_1_1__leaf_net664;
 wire clknet_0_net663;
 wire clknet_1_0__leaf_net663;
 wire clknet_1_1__leaf_net663;
 wire clknet_0_net764;
 wire clknet_1_0__leaf_net764;
 wire clknet_1_1__leaf_net764;
 wire clknet_0_net750;
 wire clknet_1_0__leaf_net750;
 wire clknet_1_1__leaf_net750;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;

 sky130_fd_sc_hd__and2_2 c100 (.A(net31),
    .B(net35),
    .X(net37));
 sky130_fd_sc_hd__and2_2 c101 (.A(net728),
    .B(net29),
    .X(net789));
 sky130_fd_sc_hd__and3_1 c102 (.A(net27),
    .B(net31),
    .C(net25),
    .X(net38));
 sky130_fd_sc_hd__and2_1 c103 (.A(net38),
    .B(net789),
    .X(net39));
 sky130_fd_sc_hd__and2_1 c104 (.A(net36),
    .B(net30),
    .X(net40));
 sky130_fd_sc_hd__and3_1 c105 (.A(net34),
    .B(net35),
    .C(net39),
    .X(net41));
 sky130_fd_sc_hd__and2_1 c106 (.A(net30),
    .B(net34),
    .X(net42));
 sky130_fd_sc_hd__and2_1 c107 (.A(net40),
    .B(net29),
    .X(net43));
 sky130_fd_sc_hd__and3_1 c108 (.A(net35),
    .B(net43),
    .C(net38),
    .X(net44));
 sky130_fd_sc_hd__a2111o_2 c109 (.A1(net44),
    .A2(net41),
    .B1(net43),
    .C1(net2),
    .D1(net33),
    .X(net45));
 sky130_fd_sc_hd__and2_0 c110 (.A(net723),
    .B(net726),
    .X(net46));
 sky130_fd_sc_hd__and2_0 c111 (.A(net46),
    .B(net724),
    .X(net774));
 sky130_fd_sc_hd__and2_0 c112 (.A(net46),
    .B(net726),
    .X(net47));
 sky130_fd_sc_hd__and2_0 c113 (.A(net721),
    .B(net32),
    .X(net48));
 sky130_fd_sc_hd__and2_0 c114 (.A(net6),
    .B(net721),
    .X(net49));
 sky130_fd_sc_hd__and2_0 c115 (.A(net30),
    .B(net46),
    .X(net50));
 sky130_fd_sc_hd__and2_0 c116 (.A(net726),
    .B(net32),
    .X(net51));
 sky130_fd_sc_hd__and2_1 c117 (.A(net49),
    .B(net5),
    .X(net52));
 sky130_fd_sc_hd__and2_2 c118 (.A(net48),
    .B(net52),
    .X(net768));
 sky130_fd_sc_hd__and2_0 c119 (.A(net32),
    .B(net52),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c120 (.A(net7),
    .B(net32),
    .X(net54));
 sky130_fd_sc_hd__and2_0 c121 (.A(net51),
    .B(net54),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c122 (.A(net47),
    .B(net54),
    .C(net768),
    .X(net56));
 sky130_fd_sc_hd__and2_0 c123 (.A(net50),
    .B(net47),
    .X(net57));
 sky130_fd_sc_hd__and2_0 c124 (.A(net47),
    .B(net768),
    .X(net751));
 sky130_fd_sc_hd__and2_0 c125 (.A(net55),
    .B(net724),
    .X(net58));
 sky130_fd_sc_hd__and2_0 c126 (.A(net54),
    .B(net58),
    .X(net59));
 sky130_fd_sc_hd__and2_0 c127 (.A(net52),
    .B(net53),
    .X(net60));
 sky130_fd_sc_hd__and2_0 c128 (.A(net53),
    .B(net58),
    .X(net61));
 sky130_fd_sc_hd__and3_1 c129 (.A(net60),
    .B(net726),
    .C(net718),
    .X(net62));
 sky130_fd_sc_hd__and2_0 c130 (.A(net56),
    .B(net52),
    .X(net63));
 sky130_fd_sc_hd__and3_1 c131 (.A(net61),
    .B(net60),
    .C(net56),
    .X(net778));
 sky130_fd_sc_hd__and2_4 c132 (.A(net686),
    .B(net676),
    .X(net64));
 sky130_fd_sc_hd__and2_0 c133 (.A(net680),
    .B(net675),
    .X(net65));
 sky130_fd_sc_hd__and2_4 c134 (.A(net683),
    .B(net729),
    .X(net66));
 sky130_fd_sc_hd__and2_4 c135 (.A(net733),
    .B(net64),
    .X(net67));
 sky130_fd_sc_hd__and2_1 c136 (.A(net676),
    .B(net680),
    .X(net68));
 sky130_fd_sc_hd__and2_4 c137 (.A(net66),
    .B(net678),
    .X(net69));
 sky130_fd_sc_hd__and2_1 c138 (.A(net732),
    .B(net67),
    .X(net70));
 sky130_fd_sc_hd__and3_4 c139 (.A(net683),
    .B(net617),
    .C(net681),
    .X(net71));
 sky130_fd_sc_hd__and2_1 c140 (.A(net71),
    .B(net66),
    .X(net72));
 sky130_fd_sc_hd__and3_4 c141 (.A(net69),
    .B(net67),
    .C(net71),
    .X(net73));
 sky130_fd_sc_hd__and2_4 c142 (.A(net69),
    .B(net73),
    .X(net74));
 sky130_fd_sc_hd__and3_1 c143 (.A(net74),
    .B(net70),
    .C(net72),
    .X(net75));
 sky130_fd_sc_hd__and2_1 c144 (.A(net68),
    .B(net72),
    .X(net76));
 sky130_fd_sc_hd__and3_4 c145 (.A(net679),
    .B(net76),
    .C(net829),
    .X(net77));
 sky130_fd_sc_hd__and3_4 c146 (.A(net66),
    .B(net75),
    .C(net69),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c147 (.A(net75),
    .B(net687),
    .C(net71),
    .X(net79));
 sky130_fd_sc_hd__or4bb_4 c148 (.A(net684),
    .B(net79),
    .C_N(net65),
    .D_N(net71),
    .X(net80));
 sky130_fd_sc_hd__and3_2 c149 (.A(net78),
    .B(net73),
    .C(net72),
    .X(net81));
 sky130_fd_sc_hd__and2_0 c150 (.A(net76),
    .B(net74),
    .X(net82));
 sky130_fd_sc_hd__and3_1 c151 (.A(net80),
    .B(net78),
    .C(net76),
    .X(net83));
 sky130_fd_sc_hd__and3_4 c152 (.A(net78),
    .B(net80),
    .C(net66),
    .X(net84));
 sky130_fd_sc_hd__a2111o_1 c153 (.A1(net83),
    .A2(net70),
    .B1(net82),
    .C1(net81),
    .D1(net74),
    .X(net85));
 sky130_fd_sc_hd__and2_0 c154 (.A(net687),
    .B(net81),
    .X(net86));
 sky130_fd_sc_hd__and2_1 c155 (.A(net696),
    .B(net81),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c156 (.A(net698),
    .B(net74),
    .X(net88));
 sky130_fd_sc_hd__and2_1 c157 (.A(net692),
    .B(net617),
    .X(net89));
 sky130_fd_sc_hd__and2_1 c158 (.A(net689),
    .B(net678),
    .X(net90));
 sky130_fd_sc_hd__and2_0 c159 (.A(net703),
    .B(net64),
    .X(net91));
 sky130_fd_sc_hd__and2_1 c160 (.A(net709),
    .B(net68),
    .X(net92));
 sky130_fd_sc_hd__and2_2 c161 (.A(net695),
    .B(net88),
    .X(net93));
 sky130_fd_sc_hd__and2_1 c162 (.A(net697),
    .B(net91),
    .X(net94));
 sky130_fd_sc_hd__and2_4 c163 (.A(net701),
    .B(net93),
    .X(net95));
 sky130_fd_sc_hd__and2_1 c164 (.A(net682),
    .B(net94),
    .X(net96));
 sky130_fd_sc_hd__and2_1 c165 (.A(net86),
    .B(net705),
    .X(net97));
 sky130_fd_sc_hd__and2_1 c166 (.A(net699),
    .B(net96),
    .X(net98));
 sky130_fd_sc_hd__and2_0 c167 (.A(net733),
    .B(net97),
    .X(net99));
 sky130_fd_sc_hd__and3_1 c168 (.A(net710),
    .B(net688),
    .C(net95),
    .X(net100));
 sky130_fd_sc_hd__and2_0 c169 (.A(net681),
    .B(net88),
    .X(net101));
 sky130_fd_sc_hd__and2_1 c170 (.A(net101),
    .B(net96),
    .X(net102));
 sky130_fd_sc_hd__and2_4 c171 (.A(net95),
    .B(net102),
    .X(net770));
 sky130_fd_sc_hd__and2_1 c172 (.A(net99),
    .B(net100),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net96),
    .A1(net770),
    .A2(net74),
    .A3(net102),
    .S0(net95),
    .S1(net92),
    .X(net104));
 sky130_fd_sc_hd__and3_2 c174 (.A(net94),
    .B(net685),
    .C(net104),
    .X(net782));
 sky130_fd_sc_hd__and2_0 c175 (.A(net87),
    .B(net102),
    .X(net105));
 sky130_fd_sc_hd__and2_1 c176 (.A(net3),
    .B(net721),
    .X(net106));
 sky130_fd_sc_hd__and2_1 c177 (.A(net79),
    .B(net705),
    .X(net107));
 sky130_fd_sc_hd__and2_0 c178 (.A(net714),
    .B(net97),
    .X(net108));
 sky130_fd_sc_hd__and2_2 c179 (.A(net74),
    .B(net714),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c180 (.A(net727),
    .B(net0),
    .X(net110));
 sky130_fd_sc_hd__and2_2 c181 (.A(net716),
    .B(net722),
    .X(net767));
 sky130_fd_sc_hd__and3_1 c182 (.A(net730),
    .B(net110),
    .C(net106),
    .X(net111));
 sky130_fd_sc_hd__and2_1 c183 (.A(net111),
    .B(net767),
    .X(net112));
 sky130_fd_sc_hd__and2_0 c184 (.A(net112),
    .B(net3),
    .X(net113));
 sky130_fd_sc_hd__and2_1 c185 (.A(net107),
    .B(net717),
    .X(net114));
 sky130_fd_sc_hd__and3_2 c186 (.A(net0),
    .B(net106),
    .C(net713),
    .X(net115));
 sky130_fd_sc_hd__and2_0 c187 (.A(net91),
    .B(net113),
    .X(net116));
 sky130_fd_sc_hd__and2_1 c188 (.A(net711),
    .B(net110),
    .X(net117));
 sky130_fd_sc_hd__and3_2 c189 (.A(net111),
    .B(net711),
    .C(net727),
    .X(net790));
 sky130_fd_sc_hd__and2_0 c190 (.A(net109),
    .B(net115),
    .X(net118));
 sky130_fd_sc_hd__and2_0 c191 (.A(net113),
    .B(net716),
    .X(net119));
 sky130_fd_sc_hd__and2_1 c192 (.A(net118),
    .B(net767),
    .X(net120));
 sky130_fd_sc_hd__and3_1 c193 (.A(net92),
    .B(net115),
    .C(net705),
    .X(net121));
 sky130_fd_sc_hd__and2_1 c194 (.A(net114),
    .B(net117),
    .X(net122));
 sky130_fd_sc_hd__and3_2 c195 (.A(net108),
    .B(net730),
    .C(net118),
    .X(net123));
 sky130_fd_sc_hd__or4bb_4 c196 (.A(net116),
    .B(net123),
    .C_N(net110),
    .D_N(net101),
    .X(net124));
 sky130_fd_sc_hd__a2111o_4 c197 (.A1(net117),
    .A2(net120),
    .B1(net724),
    .C1(net114),
    .D1(net109),
    .X(net791));
 sky130_fd_sc_hd__and2_1 c198 (.A(net688),
    .B(net791),
    .X(net125));
 sky130_fd_sc_hd__and2_0 c199 (.A(net107),
    .B(net802),
    .X(net126));
 sky130_fd_sc_hd__and2_1 c200 (.A(net829),
    .B(net123),
    .X(net127));
 sky130_fd_sc_hd__and2_0 c201 (.A(net126),
    .B(net124),
    .X(net128));
 sky130_fd_sc_hd__and2_0 c202 (.A(net731),
    .B(net127),
    .X(net129));
 sky130_fd_sc_hd__and2_1 c203 (.A(net129),
    .B(net126),
    .X(net130));
 sky130_fd_sc_hd__and2_0 c204 (.A(net119),
    .B(net73),
    .X(net131));
 sky130_fd_sc_hd__or4bb_4 c205 (.A(net90),
    .B(net24),
    .C_N(net131),
    .D_N(net88),
    .X(net132));
 sky130_fd_sc_hd__and2_1 c206 (.A(net720),
    .B(net688),
    .X(net133));
 sky130_fd_sc_hd__and2_2 c207 (.A(net88),
    .B(net130),
    .X(net741));
 sky130_fd_sc_hd__and2_1 c208 (.A(net127),
    .B(net128),
    .X(net763));
 sky130_fd_sc_hd__and2_4 c209 (.A(net132),
    .B(net16),
    .X(net134));
 sky130_fd_sc_hd__and2_0 c210 (.A(net122),
    .B(net24),
    .X(net135));
 sky130_fd_sc_hd__and2_1 c211 (.A(net4),
    .B(net135),
    .X(net775));
 sky130_fd_sc_hd__and2_1 c212 (.A(net131),
    .B(net16),
    .X(net136));
 sky130_fd_sc_hd__sdfbbn_1 c213 (.CLK_N(clknet_4_8_0_clk),
    .D(net133),
    .RESET_B(net132),
    .SCD(net741),
    .SCE(net129),
    .SET_B(net115),
    .Q(net138),
    .Q_N(net137));
 sky130_fd_sc_hd__and2_1 c214 (.A(net90),
    .B(net775),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c215 (.A(net128),
    .B(net8),
    .C(net137),
    .X(net140));
 sky130_fd_sc_hd__a2111o_2 c216 (.A1(net140),
    .A2(net139),
    .B1(net136),
    .C1(net138),
    .D1(net133),
    .X(net141));
 sky130_fd_sc_hd__dfbbn_1 c217 (.CLK_N(clknet_4_8_0_clk),
    .D(net705),
    .RESET_B(net139),
    .SET_B(net141),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__a2111o_1 c218 (.A1(net143),
    .A2(net133),
    .B1(net122),
    .C1(net15),
    .D1(net724),
    .X(net144));
 sky130_fd_sc_hd__and3_2 c219 (.A(net144),
    .B(net140),
    .C(net142),
    .X(net769));
 sky130_fd_sc_hd__and2_1 c220 (.A(net134),
    .B(net804),
    .X(net145));
 sky130_fd_sc_hd__and2_0 c221 (.A(net700),
    .B(net145),
    .X(net146));
 sky130_fd_sc_hd__and2_0 c222 (.A(net734),
    .B(net33),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net622),
    .X(net148));
 sky130_fd_sc_hd__dfbbn_1 c224 (.CLK_N(clknet_4_8_0_clk),
    .D(net722),
    .RESET_B(net146),
    .SET_B(net42),
    .Q(net149));
 sky130_fd_sc_hd__and2_1 c225 (.A(net712),
    .B(net770),
    .X(net150));
 sky130_fd_sc_hd__and2_0 c226 (.A(net145),
    .B(net790),
    .X(net151));
 sky130_fd_sc_hd__or4bb_1 c227 (.A(net855),
    .B(net804),
    .C_N(net123),
    .D_N(net125),
    .X(net152));
 sky130_fd_sc_hd__or4bb_1 c228 (.A(net40),
    .B(net87),
    .C_N(net148),
    .D_N(net37),
    .X(net153));
 sky130_fd_sc_hd__and3_1 c229 (.A(net147),
    .B(net150),
    .C(net39),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 c230 (.A(net623),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c231 (.A(net155),
    .B(net40),
    .C(net153),
    .X(net156));
 sky130_fd_sc_hd__and2_4 c232 (.A(net135),
    .B(net16),
    .X(net157));
 sky130_fd_sc_hd__and3_1 c233 (.A(net804),
    .B(net138),
    .C(net157),
    .X(net785));
 sky130_fd_sc_hd__and3_1 c234 (.A(net157),
    .B(net875),
    .C(net153),
    .X(net158));
 sky130_fd_sc_hd__a2111o_4 c235 (.A1(net156),
    .A2(net157),
    .B1(net158),
    .C1(net137),
    .D1(net134),
    .X(net159));
 sky130_fd_sc_hd__or4bb_2 c236 (.A(net41),
    .B(net145),
    .C_N(net136),
    .D_N(net157),
    .X(net160));
 sky130_fd_sc_hd__dfbbp_1 c237 (.CLK(clknet_4_10_0_clk),
    .D(net151),
    .RESET_B(net157),
    .SET_B(net160),
    .Q(net162),
    .Q_N(net161));
 sky130_fd_sc_hd__sdfxbp_1 c238 (.CLK(clknet_4_10_0_clk),
    .D(net43),
    .SCD(net852),
    .SCE(net769),
    .Q(net163));
 sky130_fd_sc_hd__sdfxbp_1 c239 (.CLK(clknet_4_10_0_clk),
    .D(net162),
    .SCD(net157),
    .SCE(net819),
    .Q(net164));
 sky130_fd_sc_hd__and3_1 c240 (.A(net163),
    .B(net162),
    .C(net157),
    .X(net788));
 sky130_fd_sc_hd__and3_1 c241 (.A(net863),
    .B(net791),
    .C(net790),
    .X(net165));
 sky130_fd_sc_hd__and2_1 c242 (.A(net63),
    .B(net36),
    .X(net166));
 sky130_fd_sc_hd__and2_0 c243 (.A(net62),
    .B(net37),
    .X(net167));
 sky130_fd_sc_hd__and2_0 c244 (.A(net16),
    .B(net708),
    .X(net168));
 sky130_fd_sc_hd__and2_1 c245 (.A(net123),
    .B(net768),
    .X(net169));
 sky130_fd_sc_hd__and2_2 c246 (.A(net35),
    .B(net169),
    .X(net777));
 sky130_fd_sc_hd__and2_1 c247 (.A(net152),
    .B(net158),
    .X(net754));
 sky130_fd_sc_hd__and2_0 c248 (.A(net37),
    .B(net777),
    .X(net170));
 sky130_fd_sc_hd__and2_0 c249 (.A(net59),
    .B(net36),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_1 c250 (.A(net627),
    .X(net762));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net158),
    .A1(net708),
    .A2(net768),
    .A3(net704),
    .S0(net724),
    .S1(net37),
    .X(net171));
 sky130_fd_sc_hd__and2_1 c252 (.A(net167),
    .B(net788),
    .X(net761));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net702),
    .A1(net36),
    .A2(net777),
    .A3(net37),
    .S0(net768),
    .S1(net154),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 c254 (.A(net627),
    .X(net173));
 sky130_fd_sc_hd__and2_0 c255 (.A(net138),
    .B(net777),
    .X(net174));
 sky130_fd_sc_hd__and2_0 c256 (.A(net172),
    .B(net37),
    .X(net783));
 sky130_fd_sc_hd__and2_1 c257 (.A(net174),
    .B(net782),
    .X(net786));
 sky130_fd_sc_hd__and2_0 c258 (.A(net168),
    .B(net777),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c259 (.A(net175),
    .B(net140),
    .C(net169),
    .X(net176));
 sky130_fd_sc_hd__buf_1 c260 (.A(net641),
    .X(net177));
 sky130_fd_sc_hd__and2_1 c261 (.A(net177),
    .B(net52),
    .X(net757));
 sky130_fd_sc_hd__sdfbbn_1 c262 (.CLK_N(clknet_4_10_0_clk),
    .D(net173),
    .RESET_B(net177),
    .SCD(net757),
    .SCE(net777),
    .SET_B(net786),
    .Q(net780),
    .Q_N(net178));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net170),
    .A1(net178),
    .A2(net169),
    .A3(net786),
    .S0(net777),
    .S1(net52),
    .X(net179));
 sky130_fd_sc_hd__and2_1 c264 (.A(net82),
    .B(net76),
    .X(net180));
 sky130_fd_sc_hd__and2_4 c265 (.A(net65),
    .B(net84),
    .X(net181));
 sky130_fd_sc_hd__and2_1 c266 (.A(net69),
    .B(net82),
    .X(net182));
 sky130_fd_sc_hd__and2_1 c267 (.A(net180),
    .B(net674),
    .X(net183));
 sky130_fd_sc_hd__and2_4 c268 (.A(net80),
    .B(net71),
    .X(net184));
 sky130_fd_sc_hd__and2_2 c269 (.A(net184),
    .B(net182),
    .X(net185));
 sky130_fd_sc_hd__and2_2 c270 (.A(net732),
    .B(net729),
    .X(net772));
 sky130_fd_sc_hd__and2_1 c271 (.A(net181),
    .B(net85),
    .X(net186));
 sky130_fd_sc_hd__and2_1 c272 (.A(net707),
    .B(net71),
    .X(net187));
 sky130_fd_sc_hd__and2_1 c273 (.A(net707),
    .B(net71),
    .X(net188));
 sky130_fd_sc_hd__and2_0 c274 (.A(net186),
    .B(net64),
    .X(net189));
 sky130_fd_sc_hd__and3_1 c275 (.A(net186),
    .B(net183),
    .C(net181),
    .X(net190));
 sky130_fd_sc_hd__and2_1 c276 (.A(net190),
    .B(net188),
    .X(net191));
 sky130_fd_sc_hd__or4bb_4 c277 (.A(net188),
    .B(net617),
    .C_N(net187),
    .D_N(net794),
    .X(net192));
 sky130_fd_sc_hd__and3_1 c278 (.A(net191),
    .B(net73),
    .C(net794),
    .X(net193));
 sky130_fd_sc_hd__and2_0 c279 (.A(net71),
    .B(net183),
    .X(net194));
 sky130_fd_sc_hd__and2_1 c280 (.A(net189),
    .B(net184),
    .X(net195));
 sky130_fd_sc_hd__and2_1 c281 (.A(net186),
    .B(net190),
    .X(net196));
 sky130_fd_sc_hd__and2_1 c282 (.A(net195),
    .B(net187),
    .X(net197));
 sky130_fd_sc_hd__and3_1 c283 (.A(net85),
    .B(net194),
    .C(net192),
    .X(net198));
 sky130_fd_sc_hd__and2_2 c284 (.A(net198),
    .B(net69),
    .X(net199));
 sky130_fd_sc_hd__or4bb_4 c285 (.A(net197),
    .B(net190),
    .C_N(net794),
    .D_N(net186),
    .X(net200));
 sky130_fd_sc_hd__and2_1 c286 (.A(net617),
    .B(net182),
    .X(net201));
 sky130_fd_sc_hd__and3_1 c287 (.A(net182),
    .B(net96),
    .C(net201),
    .X(net202));
 sky130_fd_sc_hd__and2_0 c288 (.A(net190),
    .B(net685),
    .X(net203));
 sky130_fd_sc_hd__and2_0 c289 (.A(net68),
    .B(net702),
    .X(net204));
 sky130_fd_sc_hd__and2_1 c290 (.A(net197),
    .B(net95),
    .X(net205));
 sky130_fd_sc_hd__and2_4 c291 (.A(net189),
    .B(net192),
    .X(net206));
 sky130_fd_sc_hd__and3_1 c292 (.A(net202),
    .B(net98),
    .C(net205),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c293 (.A(net690),
    .B(net199),
    .X(net744));
 sky130_fd_sc_hd__and2_0 c294 (.A(net203),
    .B(net188),
    .X(net208));
 sky130_fd_sc_hd__buf_2 c295 (.A(net671),
    .X(net746));
 sky130_fd_sc_hd__and3_1 c296 (.A(net199),
    .B(net78),
    .C(net192),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c297 (.A(net94),
    .B(net782),
    .C(net206),
    .X(net210));
 sky130_fd_sc_hd__and3_4 c298 (.A(net194),
    .B(net185),
    .C(net794),
    .X(net211));
 sky130_fd_sc_hd__and2_0 c299 (.A(net691),
    .B(net209),
    .X(net212));
 sky130_fd_sc_hd__and2_1 c300 (.A(net676),
    .B(net206),
    .X(net213));
 sky130_fd_sc_hd__and2_2 c301 (.A(net86),
    .B(net820),
    .X(net214));
 sky130_fd_sc_hd__sdfbbp_1 c302 (.CLK(clknet_4_0_0_clk),
    .D(net211),
    .RESET_B(net204),
    .SCD(net214),
    .SCE(net213),
    .SET_B(net206),
    .Q(net216),
    .Q_N(net215));
 sky130_fd_sc_hd__and3_1 c303 (.A(net64),
    .B(net216),
    .C(net211),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 c304 (.A(net671),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c305 (.A(net675),
    .B(net217),
    .C(net95),
    .X(net219));
 sky130_fd_sc_hd__a2111o_4 c306 (.A1(net204),
    .A2(net94),
    .B1(net64),
    .C1(net219),
    .D1(net206),
    .X(net220));
 sky130_fd_sc_hd__a2111o_4 c307 (.A1(net205),
    .A2(net217),
    .B1(net103),
    .C1(net215),
    .D1(net219),
    .X(net221));
 sky130_fd_sc_hd__and2_1 c308 (.A(net102),
    .B(net208),
    .X(net222));
 sky130_fd_sc_hd__and2_0 c309 (.A(net105),
    .B(net872),
    .X(net223));
 sky130_fd_sc_hd__and2_1 c310 (.A(net208),
    .B(net124),
    .X(net224));
 sky130_fd_sc_hd__and2_0 c311 (.A(net188),
    .B(net2),
    .X(net225));
 sky130_fd_sc_hd__and2_0 c312 (.A(net686),
    .B(net224),
    .X(net226));
 sky130_fd_sc_hd__and2_1 c313 (.A(net216),
    .B(net220),
    .X(net227));
 sky130_fd_sc_hd__and3_1 c314 (.A(net685),
    .B(net734),
    .C(net746),
    .X(net228));
 sky130_fd_sc_hd__and3_4 c315 (.A(net103),
    .B(net215),
    .C(net89),
    .X(net776));
 sky130_fd_sc_hd__sdfxtp_1 c316 (.CLK(clknet_4_2_0_clk),
    .D(net226),
    .SCD(net678),
    .SCE(net216),
    .Q(net229));
 sky130_fd_sc_hd__and2_0 c317 (.A(net228),
    .B(net227),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c318 (.A(net227),
    .B(net821),
    .X(net231));
 sky130_fd_sc_hd__buf_1 c319 (.A(net613),
    .X(net232));
 sky130_fd_sc_hd__buf_1 c320 (.A(net612),
    .X(net233));
 sky130_fd_sc_hd__sdfxtp_1 c321 (.CLK(clknet_4_2_0_clk),
    .D(net228),
    .SCD(net226),
    .SCE(net223),
    .Q(net234));
 sky130_fd_sc_hd__sdfxtp_1 c322 (.CLK(clknet_4_2_0_clk),
    .D(net230),
    .SCD(net866),
    .SCE(net721),
    .Q(net235));
 sky130_fd_sc_hd__and3_2 c323 (.A(net223),
    .B(net235),
    .C(net232),
    .X(net236));
 sky130_fd_sc_hd__dfbbn_1 c324 (.CLK_N(clknet_4_2_0_clk),
    .D(net225),
    .RESET_B(net235),
    .SET_B(net231),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__a2111o_1 c325 (.A1(net233),
    .A2(net236),
    .B1(net717),
    .C1(net229),
    .D1(net776),
    .X(net239));
 sky130_fd_sc_hd__and3_1 c326 (.A(net868),
    .B(net239),
    .C(net225),
    .X(net240));
 sky130_fd_sc_hd__and3_1 c327 (.A(net120),
    .B(net240),
    .C(net105),
    .X(net241));
 sky130_fd_sc_hd__dfbbn_1 c328 (.CLK_N(clknet_4_8_0_clk),
    .D(net241),
    .RESET_B(net239),
    .SET_B(net233),
    .Q(net243),
    .Q_N(net242));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net232),
    .A1(net240),
    .A2(net236),
    .A3(net242),
    .S0(net241),
    .S1(net124),
    .X(net244));
 sky130_fd_sc_hd__and2_0 c330 (.A(net229),
    .B(net227),
    .X(net245));
 sky130_fd_sc_hd__and2_1 c331 (.A(net678),
    .B(net243),
    .X(net246));
 sky130_fd_sc_hd__and3_2 c332 (.A(net246),
    .B(net763),
    .C(net115),
    .X(net743));
 sky130_fd_sc_hd__and2_0 c333 (.A(net729),
    .B(net240),
    .X(net247));
 sky130_fd_sc_hd__a2111o_1 c334 (.A1(net124),
    .A2(net775),
    .B1(net109),
    .C1(net133),
    .D1(net794),
    .X(net248));
 sky130_fd_sc_hd__and2_0 c335 (.A(net144),
    .B(net229),
    .X(net249));
 sky130_fd_sc_hd__and3_1 c336 (.A(net181),
    .B(net106),
    .C(net15),
    .X(net250));
 sky130_fd_sc_hd__and3_2 c337 (.A(net249),
    .B(net239),
    .C(net248),
    .X(net735));
 sky130_fd_sc_hd__dfbbp_1 c338 (.CLK(clknet_4_8_0_clk),
    .D(net245),
    .RESET_B(net106),
    .SET_B(net246),
    .Q(net251));
 sky130_fd_sc_hd__and2_1 c339 (.A(net239),
    .B(net78),
    .X(net252));
 sky130_fd_sc_hd__and2_1 c340 (.A(net78),
    .B(net763),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 c341 (.A(net624),
    .X(net253));
 sky130_fd_sc_hd__and2_0 c342 (.A(net252),
    .B(net729),
    .X(net254));
 sky130_fd_sc_hd__and3_1 c343 (.A(net115),
    .B(net725),
    .C(net229),
    .X(net255));
 sky130_fd_sc_hd__and2_1 c344 (.A(net240),
    .B(net248),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c345 (.A(net250),
    .B(net678),
    .C(net734),
    .X(net257));
 sky130_fd_sc_hd__and2_0 c346 (.A(net255),
    .B(net252),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net624),
    .X(net259));
 sky130_fd_sc_hd__and2_0 c348 (.A(net257),
    .B(net645),
    .X(net260));
 sky130_fd_sc_hd__sdfxbp_2 c349 (.CLK(clknet_4_8_0_clk),
    .D(net260),
    .SCD(net227),
    .SCE(net245),
    .Q(net262),
    .Q_N(net261));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net258),
    .A1(net130),
    .A2(net257),
    .A3(net260),
    .S0(net261),
    .S1(net246),
    .X(net263));
 sky130_fd_sc_hd__sdfxbp_1 c351 (.CLK(clknet_4_12_0_clk),
    .D(net254),
    .SCD(net247),
    .SCE(net854),
    .Q(net265),
    .Q_N(net264));
 sky130_fd_sc_hd__and2_4 c352 (.A(net153),
    .B(net261),
    .X(net266));
 sky130_fd_sc_hd__and2_0 c353 (.A(net150),
    .B(net77),
    .X(net267));
 sky130_fd_sc_hd__and2_1 c354 (.A(net873),
    .B(net259),
    .X(net755));
 sky130_fd_sc_hd__and2_0 c355 (.A(net33),
    .B(net721),
    .X(net268));
 sky130_fd_sc_hd__buf_1 c356 (.A(net629),
    .X(net269));
 sky130_fd_sc_hd__and2_1 c357 (.A(net136),
    .B(net872),
    .X(net270));
 sky130_fd_sc_hd__and2_2 c358 (.A(net42),
    .B(net125),
    .X(net271));
 sky130_fd_sc_hd__and2_0 c359 (.A(net268),
    .B(net718),
    .X(net272));
 sky130_fd_sc_hd__and2_0 c360 (.A(net234),
    .B(net270),
    .X(net273));
 sky130_fd_sc_hd__sdfrbp_1 c361 (.CLK(clknet_4_10_0_clk),
    .D(net165),
    .RESET_B(net734),
    .SCD(net271),
    .SCE(net160),
    .Q(net275),
    .Q_N(net274));
 sky130_fd_sc_hd__and2_0 c362 (.A(net272),
    .B(net262),
    .X(net276));
 sky130_fd_sc_hd__and3_2 c363 (.A(net130),
    .B(net834),
    .C(net271),
    .X(net765));
 sky130_fd_sc_hd__and2_0 c364 (.A(net273),
    .B(net795),
    .X(net277));
 sky130_fd_sc_hd__buf_1 c365 (.A(net629),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 c366 (.A(net641),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net106),
    .A1(net755),
    .A2(net276),
    .A3(net150),
    .S0(net271),
    .S1(net769),
    .X(net280));
 sky130_fd_sc_hd__and2_1 c368 (.A(net277),
    .B(net278),
    .X(net781));
 sky130_fd_sc_hd__and3_1 c369 (.A(net276),
    .B(net873),
    .C(net795),
    .X(net281));
 sky130_fd_sc_hd__dfrbp_1 c370 (.CLK(clknet_4_11_0_clk),
    .D(net281),
    .RESET_B(net765),
    .Q(net283),
    .Q_N(net282));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net874),
    .A1(net275),
    .A2(net281),
    .A3(net234),
    .S0(net271),
    .S1(net647),
    .X(net284));
 sky130_fd_sc_hd__and2_1 c372 (.A(net284),
    .B(net271),
    .X(net771));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net279),
    .A1(net281),
    .A2(net743),
    .A3(net781),
    .S0(net282),
    .S1(net860),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net57),
    .A1(net177),
    .A2(net786),
    .A3(net828),
    .S0(net741),
    .S1(net761),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net154),
    .A1(net77),
    .A2(net765),
    .A3(net767),
    .S0(net177),
    .S1(clknet_1_0__leaf_net750),
    .X(net287));
 sky130_fd_sc_hd__sdfbbn_1 c394 (.CLK_N(clknet_4_10_0_clk),
    .D(net166),
    .RESET_B(net721),
    .SCD(net754),
    .SCE(clknet_1_0__leaf_net750),
    .SET_B(clknet_1_0__leaf_net764),
    .Q(net784),
    .Q_N(net288));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net267),
    .A1(net791),
    .A2(net288),
    .A3(net757),
    .S0(clknet_1_1__leaf_net750),
    .S1(clknet_1_0__leaf_net764),
    .X(net787));
 sky130_fd_sc_hd__and2_0 c396 (.A(net198),
    .B(net81),
    .X(net289));
 sky130_fd_sc_hd__and2_0 c397 (.A(net684),
    .B(net183),
    .X(net290));
 sky130_fd_sc_hd__and2_0 c398 (.A(net289),
    .B(net729),
    .X(net291));
 sky130_fd_sc_hd__and2_1 c399 (.A(net289),
    .B(net70),
    .X(net292));
 sky130_fd_sc_hd__and2_4 c400 (.A(net200),
    .B(net290),
    .X(net293));
 sky130_fd_sc_hd__and2_1 c401 (.A(net292),
    .B(net193),
    .X(net294));
 sky130_fd_sc_hd__and2_1 c402 (.A(net76),
    .B(net294),
    .X(net295));
 sky130_fd_sc_hd__and2_0 c403 (.A(net291),
    .B(net81),
    .X(net296));
 sky130_fd_sc_hd__and2_4 c404 (.A(net187),
    .B(net184),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c405 (.A(net183),
    .B(net292),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 c406 (.A(net611),
    .X(net299));
 sky130_fd_sc_hd__and2_4 c407 (.A(net296),
    .B(net298),
    .X(net300));
 sky130_fd_sc_hd__and2_2 c408 (.A(net292),
    .B(net187),
    .X(net301));
 sky130_fd_sc_hd__and2_2 c409 (.A(net294),
    .B(net300),
    .X(net302));
 sky130_fd_sc_hd__and2_1 c410 (.A(net298),
    .B(net185),
    .X(net303));
 sky130_fd_sc_hd__and2_1 c411 (.A(net301),
    .B(net303),
    .X(net304));
 sky130_fd_sc_hd__dlymetal6s2s_1 c412 (.A(net611),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 c413 (.A(net639),
    .X(net306));
 sky130_fd_sc_hd__and3_1 c414 (.A(net305),
    .B(net291),
    .C(net306),
    .X(net307));
 sky130_fd_sc_hd__and2_0 c415 (.A(net307),
    .B(net290),
    .X(net308));
 sky130_fd_sc_hd__and2_0 c416 (.A(net290),
    .B(net305),
    .X(net309));
 sky130_fd_sc_hd__and3_1 c417 (.A(net308),
    .B(net296),
    .C(net305),
    .X(net310));
 sky130_fd_sc_hd__sdfrbp_1 c418 (.CLK(clknet_4_0_0_clk),
    .D(net309),
    .RESET_B(net303),
    .SCD(net310),
    .SCE(net95),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__and2_2 c419 (.A(net218),
    .B(net201),
    .X(net313));
 sky130_fd_sc_hd__and3_1 c420 (.A(net312),
    .B(net95),
    .C(net301),
    .X(net314));
 sky130_fd_sc_hd__sdfxtp_1 c421 (.CLK(clknet_4_0_0_clk),
    .D(net310),
    .SCD(net81),
    .SCE(net313),
    .Q(net315));
 sky130_fd_sc_hd__and2_0 c422 (.A(net193),
    .B(net823),
    .X(net316));
 sky130_fd_sc_hd__or4bb_1 c423 (.A(net210),
    .B(net211),
    .C_N(net70),
    .D_N(net313),
    .X(net317));
 sky130_fd_sc_hd__and3_1 c424 (.A(net211),
    .B(net315),
    .C(net729),
    .X(net318));
 sky130_fd_sc_hd__and2_1 c425 (.A(net201),
    .B(net312),
    .X(net319));
 sky130_fd_sc_hd__and2_0 c426 (.A(net209),
    .B(net307),
    .X(net320));
 sky130_fd_sc_hd__and2_1 c427 (.A(net320),
    .B(net193),
    .X(net321));
 sky130_fd_sc_hd__a2111o_2 c428 (.A1(net219),
    .A2(net318),
    .B1(net81),
    .C1(net311),
    .D1(net211),
    .X(net322));
 sky130_fd_sc_hd__sdfrtn_1 c429 (.CLK_N(clknet_4_0_0_clk),
    .D(net70),
    .RESET_B(net193),
    .SCD(net310),
    .SCE(net220),
    .Q(net323));
 sky130_fd_sc_hd__and3_1 c430 (.A(net306),
    .B(net313),
    .C(net210),
    .X(net324));
 sky130_fd_sc_hd__and2_1 c431 (.A(net299),
    .B(net324),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net314),
    .A1(net303),
    .A2(net320),
    .A3(net325),
    .S0(net321),
    .S1(net211),
    .X(net326));
 sky130_fd_sc_hd__and2_1 c433 (.A(net104),
    .B(net201),
    .X(net327));
 sky130_fd_sc_hd__sdfrtp_1 c434 (.CLK(clknet_4_1_0_clk),
    .D(net317),
    .RESET_B(net323),
    .SCD(net302),
    .SCE(net792),
    .Q(net328));
 sky130_fd_sc_hd__buf_1 c435 (.A(net619),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net316),
    .A1(net313),
    .A2(net322),
    .A3(net325),
    .S0(net329),
    .S1(net794),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 c437 (.A(net619),
    .X(net331));
 sky130_fd_sc_hd__and3_1 c438 (.A(net331),
    .B(net313),
    .C(net792),
    .X(net332));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net323),
    .A1(net792),
    .A2(net332),
    .A3(net313),
    .S0(net794),
    .S1(net649),
    .X(net758));
 sky130_fd_sc_hd__and2_1 c440 (.A(net318),
    .B(net224),
    .X(net333));
 sky130_fd_sc_hd__and2_0 c441 (.A(net313),
    .B(net717),
    .X(net334));
 sky130_fd_sc_hd__a2111o_2 c442 (.A1(net674),
    .A2(net322),
    .B1(net222),
    .C1(net725),
    .D1(net327),
    .X(net335));
 sky130_fd_sc_hd__buf_1 c443 (.A(net642),
    .X(net336));
 sky130_fd_sc_hd__and2_4 c444 (.A(net329),
    .B(net220),
    .X(net337));
 sky130_fd_sc_hd__sdfxtp_1 c445 (.CLK(clknet_4_3_0_clk),
    .D(net336),
    .SCD(net236),
    .SCE(net221),
    .Q(net338));
 sky130_fd_sc_hd__clkbuf_1 c446 (.A(net618),
    .X(net339));
 sky130_fd_sc_hd__and3_2 c447 (.A(net110),
    .B(net236),
    .C(net725),
    .X(net340));
 sky130_fd_sc_hd__and3_1 c448 (.A(net337),
    .B(net336),
    .C(net93),
    .X(net341));
 sky130_fd_sc_hd__sdfxtp_1 c449 (.CLK(clknet_4_1_0_clk),
    .D(net335),
    .SCD(net212),
    .SCE(net715),
    .Q(net342));
 sky130_fd_sc_hd__and3_1 c450 (.A(net339),
    .B(net336),
    .C(net222),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 c451 (.A(net618),
    .X(net344));
 sky130_fd_sc_hd__and2_4 c452 (.A(net823),
    .B(net342),
    .X(net345));
 sky130_fd_sc_hd__and3_4 c453 (.A(net342),
    .B(net337),
    .C(net303),
    .X(net346));
 sky130_fd_sc_hd__dfbbn_1 c454 (.CLK_N(clknet_4_9_0_clk),
    .D(net843),
    .RESET_B(net322),
    .SET_B(net345),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__sdfbbn_1 c455 (.CLK_N(clknet_4_12_0_clk),
    .D(net341),
    .RESET_B(net839),
    .SCD(net346),
    .SCE(net776),
    .SET_B(net335),
    .Q(net350),
    .Q_N(net349));
 sky130_fd_sc_hd__buf_1 c456 (.A(net640),
    .X(net351));
 sky130_fd_sc_hd__dfbbn_1 c457 (.CLK_N(clknet_4_3_0_clk),
    .D(net212),
    .RESET_B(net93),
    .SET_B(net346),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__and3_1 c458 (.A(net222),
    .B(net352),
    .C(net347),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net303),
    .A1(net353),
    .A2(net339),
    .A3(net708),
    .S0(net333),
    .S1(net242),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net89),
    .A1(net353),
    .A2(net345),
    .A3(net236),
    .S0(net350),
    .S1(net650),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net340),
    .A1(net725),
    .A2(net341),
    .A3(net345),
    .S0(net651),
    .S1(net653),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 c462 (.A(net621),
    .X(net358));
 sky130_fd_sc_hd__and2_2 c463 (.A(net93),
    .B(net358),
    .X(net359));
 sky130_fd_sc_hd__dfbbp_1 c464 (.CLK(clknet_4_9_0_clk),
    .D(net818),
    .RESET_B(net9),
    .SET_B(net830),
    .Q(net360));
 sky130_fd_sc_hd__and2_1 c465 (.A(net253),
    .B(net351),
    .X(net361));
 sky130_fd_sc_hd__and2_2 c466 (.A(net8),
    .B(net262),
    .X(net362));
 sky130_fd_sc_hd__and3_1 c467 (.A(net857),
    .B(net704),
    .C(net674),
    .X(net363));
 sky130_fd_sc_hd__and2_1 c468 (.A(net360),
    .B(net133),
    .X(net364));
 sky130_fd_sc_hd__and2_0 c469 (.A(net364),
    .B(net746),
    .X(net365));
 sky130_fd_sc_hd__and3_1 c470 (.A(net248),
    .B(net359),
    .C(net708),
    .X(net366));
 sky130_fd_sc_hd__or4bb_4 c471 (.A(net359),
    .B(net93),
    .C_N(net185),
    .D_N(net252),
    .X(net748));
 sky130_fd_sc_hd__and2_2 c472 (.A(net363),
    .B(net364),
    .X(net760));
 sky130_fd_sc_hd__and2_2 c473 (.A(net803),
    .B(net359),
    .X(net756));
 sky130_fd_sc_hd__and3_1 c474 (.A(net139),
    .B(net790),
    .C(net2),
    .X(net367));
 sky130_fd_sc_hd__sdfrtp_1 c475 (.CLK(clknet_4_9_0_clk),
    .D(net367),
    .RESET_B(net760),
    .SCD(net364),
    .SCE(net748),
    .Q(net368));
 sky130_fd_sc_hd__sdfrtp_1 c476 (.CLK(clknet_4_9_0_clk),
    .D(net840),
    .RESET_B(net835),
    .SCD(net756),
    .SCE(net817),
    .Q(net369));
 sky130_fd_sc_hd__or4bb_1 c477 (.A(net369),
    .B(net344),
    .C_N(net756),
    .D_N(net109),
    .X(net370));
 sky130_fd_sc_hd__dlymetal6s2s_1 c478 (.A(net862),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net344),
    .A1(net2),
    .A2(net243),
    .A3(net366),
    .S0(net8),
    .S1(net300),
    .X(net372));
 sky130_fd_sc_hd__or4bb_1 c480 (.A(net364),
    .B(net359),
    .C_N(net264),
    .D_N(net655),
    .X(net373));
 sky130_fd_sc_hd__sdfxbp_1 c481 (.CLK(clknet_4_9_0_clk),
    .D(net365),
    .SCD(net366),
    .SCE(net791),
    .Q(net375),
    .Q_N(net374));
 sky130_fd_sc_hd__sdfsbp_1 c482 (.CLK(clknet_4_12_0_clk),
    .D(net373),
    .SCD(net361),
    .SCE(net359),
    .SET_B(net256),
    .Q(net376));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net376),
    .A1(net756),
    .A2(net364),
    .A3(net302),
    .S0(net362),
    .S1(net655),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 c484 (.A(net615),
    .X(net378));
 sky130_fd_sc_hd__and3_1 c485 (.A(net375),
    .B(net266),
    .C(net378),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 c486 (.A(net614),
    .X(net752));
 sky130_fd_sc_hd__and3_1 c487 (.A(net283),
    .B(net300),
    .C(net266),
    .X(net380));
 sky130_fd_sc_hd__sdfxbp_1 c488 (.CLK(clknet_4_12_0_clk),
    .D(net366),
    .SCD(net302),
    .SCE(net269),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__sdfbbp_1 c489 (.CLK(clknet_4_14_0_clk),
    .D(net845),
    .RESET_B(net865),
    .SCD(net340),
    .SCE(net346),
    .SET_B(net371),
    .Q(net384),
    .Q_N(net383));
 sky130_fd_sc_hd__and3_1 c490 (.A(net278),
    .B(net381),
    .C(net708),
    .X(net385));
 sky130_fd_sc_hd__and2_0 c491 (.A(net385),
    .B(net266),
    .X(net386));
 sky130_fd_sc_hd__sdfxtp_1 c492 (.CLK(clknet_4_11_0_clk),
    .D(net259),
    .SCD(net221),
    .SCE(net2),
    .Q(net766));
 sky130_fd_sc_hd__sdfxtp_2 c493 (.CLK(clknet_4_11_0_clk),
    .D(net39),
    .SCD(net380),
    .SCE(net385),
    .Q(net387));
 sky130_fd_sc_hd__sdfxtp_1 c494 (.CLK(clknet_4_11_0_clk),
    .D(net854),
    .SCD(net748),
    .SCE(net760),
    .Q(net388));
 sky130_fd_sc_hd__and3_1 c495 (.A(net388),
    .B(net379),
    .C(net745),
    .X(net389));
 sky130_fd_sc_hd__and3_1 c496 (.A(net389),
    .B(net278),
    .C(net388),
    .X(net753));
 sky130_fd_sc_hd__and3_2 c497 (.A(net9),
    .B(net262),
    .C(net378),
    .X(net390));
 sky130_fd_sc_hd__a2111o_1 c498 (.A1(net270),
    .A2(net388),
    .B1(net269),
    .C1(net385),
    .D1(net795),
    .X(net391));
 sky130_fd_sc_hd__and3_1 c499 (.A(net729),
    .B(net382),
    .C(net390),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net125),
    .A1(net159),
    .A2(net390),
    .A3(net378),
    .S0(net753),
    .S1(net758),
    .X(net393));
 sky130_fd_sc_hd__and3_1 c501 (.A(net391),
    .B(net379),
    .C(net383),
    .X(net394));
 sky130_fd_sc_hd__and3_1 c502 (.A(net394),
    .B(net392),
    .C(net125),
    .X(net395));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net395),
    .A1(net159),
    .A2(net753),
    .A3(net776),
    .S0(net387),
    .S1(net378),
    .X(net396));
 sky130_fd_sc_hd__and3_1 c504 (.A(net386),
    .B(net378),
    .C(net387),
    .X(net397));
 sky130_fd_sc_hd__and3_1 c505 (.A(net397),
    .B(net340),
    .C(net657),
    .X(net398));
 sky130_fd_sc_hd__buf_1 c528 (.A(net633),
    .X(net399));
 sky130_fd_sc_hd__and2_1 c529 (.A(net72),
    .B(net185),
    .X(net400));
 sky130_fd_sc_hd__and2_1 c530 (.A(net400),
    .B(net301),
    .X(net401));
 sky130_fd_sc_hd__and2_4 c531 (.A(net297),
    .B(net718),
    .X(net402));
 sky130_fd_sc_hd__and2_1 c532 (.A(net196),
    .B(net300),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 c533 (.A(net832),
    .X(net404));
 sky130_fd_sc_hd__and2_1 c534 (.A(net298),
    .B(net404),
    .X(net405));
 sky130_fd_sc_hd__dfbbn_1 c535 (.CLK_N(clknet_4_4_0_clk),
    .D(net405),
    .RESET_B(net403),
    .SET_B(net196),
    .Q(net406));
 sky130_fd_sc_hd__dfrbp_1 c536 (.CLK(clknet_4_4_0_clk),
    .D(net403),
    .RESET_B(net297),
    .Q(net407));
 sky130_fd_sc_hd__and2_0 c537 (.A(net184),
    .B(net67),
    .X(net408));
 sky130_fd_sc_hd__dfbbn_1 c538 (.CLK_N(clknet_4_1_0_clk),
    .D(net408),
    .RESET_B(net403),
    .SET_B(net297),
    .Q(net409));
 sky130_fd_sc_hd__and3_2 c539 (.A(net294),
    .B(net399),
    .C(net402),
    .X(net410));
 sky130_fd_sc_hd__dfbbp_1 c540 (.CLK(clknet_4_4_0_clk),
    .D(net406),
    .RESET_B(net304),
    .SET_B(net298),
    .Q(net742),
    .Q_N(net411));
 sky130_fd_sc_hd__sdfxbp_1 c541 (.CLK(clknet_4_4_0_clk),
    .D(net401),
    .SCD(net295),
    .SCE(net411),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__dfrtn_1 c542 (.CLK_N(clknet_4_4_0_clk),
    .D(net407),
    .RESET_B(net403),
    .Q(net414));
 sky130_fd_sc_hd__and2_1 c543 (.A(net409),
    .B(net800),
    .X(net415));
 sky130_fd_sc_hd__dfrtp_1 c544 (.CLK(clknet_4_4_0_clk),
    .D(net410),
    .RESET_B(net405),
    .Q(net416));
 sky130_fd_sc_hd__and2_0 c545 (.A(net404),
    .B(net72),
    .X(net417));
 sky130_fd_sc_hd__and2_0 c546 (.A(net864),
    .B(net415),
    .X(net418));
 sky130_fd_sc_hd__and2_1 c547 (.A(net413),
    .B(net418),
    .X(net419));
 sky130_fd_sc_hd__and3_1 c548 (.A(net412),
    .B(net400),
    .C(net418),
    .X(net420));
 sky130_fd_sc_hd__sdfxbp_1 c549 (.CLK(clknet_4_4_0_clk),
    .D(net418),
    .SCD(net410),
    .SCE(net400),
    .Q(net422),
    .Q_N(net421));
 sky130_fd_sc_hd__and2_0 c550 (.A(net324),
    .B(net307),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c551 (.A(net637),
    .X(net424));
 sky130_fd_sc_hd__and2_2 c552 (.A(net213),
    .B(net307),
    .X(net425));
 sky130_fd_sc_hd__and2_0 c553 (.A(net424),
    .B(net858),
    .X(net426));
 sky130_fd_sc_hd__and2_1 c554 (.A(net417),
    .B(net98),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net636),
    .X(net428));
 sky130_fd_sc_hd__and3_1 c556 (.A(net694),
    .B(net425),
    .C(net427),
    .X(net429));
 sky130_fd_sc_hd__dfrtp_1 c557 (.CLK(clknet_4_6_0_clk),
    .D(net321),
    .RESET_B(net425),
    .Q(net430));
 sky130_fd_sc_hd__and2_0 c558 (.A(net425),
    .B(net300),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c559 (.A(net427),
    .B(net426),
    .C(net300),
    .X(net432));
 sky130_fd_sc_hd__and2_0 c560 (.A(net693),
    .B(net300),
    .X(net433));
 sky130_fd_sc_hd__sdfxtp_1 c561 (.CLK(clknet_4_1_0_clk),
    .D(net432),
    .SCD(net425),
    .SCE(net792),
    .Q(net434));
 sky130_fd_sc_hd__and2_2 c562 (.A(net100),
    .B(net323),
    .X(net435));
 sky130_fd_sc_hd__dfrtp_1 c563 (.CLK(clknet_4_6_0_clk),
    .D(net429),
    .RESET_B(net425),
    .Q(net436));
 sky130_fd_sc_hd__and3_4 c564 (.A(net434),
    .B(net435),
    .C(net323),
    .X(net437));
 sky130_fd_sc_hd__and2_0 c565 (.A(net414),
    .B(net437),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net428),
    .A1(net433),
    .A2(net694),
    .A3(net301),
    .S0(net323),
    .S1(net425),
    .X(net439));
 sky130_fd_sc_hd__and2_0 c567 (.A(net414),
    .B(net658),
    .X(net440));
 sky130_fd_sc_hd__a2111o_1 c568 (.A1(net426),
    .A2(net437),
    .B1(net425),
    .C1(net746),
    .D1(net322),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net438),
    .A1(net425),
    .A2(net437),
    .A3(net746),
    .S0(net441),
    .S1(net323),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net401),
    .A1(net98),
    .A2(net427),
    .A3(net307),
    .S0(net435),
    .S1(net859),
    .X(net443));
 sky130_fd_sc_hd__dfsbp_1 c571 (.CLK(clknet_4_6_0_clk),
    .D(net431),
    .SET_B(net441),
    .Q(net445),
    .Q_N(net444));
 sky130_fd_sc_hd__and2_1 c572 (.A(net718),
    .B(net73),
    .X(net446));
 sky130_fd_sc_hd__and2_0 c573 (.A(net419),
    .B(net338),
    .X(net447));
 sky130_fd_sc_hd__a2111o_1 c574 (.A1(net192),
    .A2(net2),
    .B1(net419),
    .C1(net340),
    .D1(net793),
    .X(net736));
 sky130_fd_sc_hd__and3_1 c575 (.A(net742),
    .B(net436),
    .C(net653),
    .X(net448));
 sky130_fd_sc_hd__and2_0 c576 (.A(net445),
    .B(net654),
    .X(net449));
 sky130_fd_sc_hd__and2_0 c577 (.A(net338),
    .B(net436),
    .X(net450));
 sky130_fd_sc_hd__and2_1 c578 (.A(net793),
    .B(net654),
    .X(net451));
 sky130_fd_sc_hd__and3_1 c579 (.A(net449),
    .B(net192),
    .C(net793),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 c580 (.A(net631),
    .X(net453));
 sky130_fd_sc_hd__and2_1 c581 (.A(net436),
    .B(net445),
    .X(net454));
 sky130_fd_sc_hd__and2_0 c582 (.A(net452),
    .B(net870),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 c583 (.A(net631),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c584 (.A(net643),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net224),
    .A1(net448),
    .A2(net718),
    .A3(net444),
    .S0(net708),
    .S1(net345),
    .X(net458));
 sky130_fd_sc_hd__and2_1 c586 (.A(net450),
    .B(net448),
    .X(net459));
 sky130_fd_sc_hd__and3_2 c587 (.A(net453),
    .B(net459),
    .C(net454),
    .X(net740));
 sky130_fd_sc_hd__and3_1 c588 (.A(net206),
    .B(net451),
    .C(net459),
    .X(net460));
 sky130_fd_sc_hd__and3_1 c589 (.A(net220),
    .B(net459),
    .C(net451),
    .X(net461));
 sky130_fd_sc_hd__and3_1 c590 (.A(net448),
    .B(net459),
    .C(net740),
    .X(net462));
 sky130_fd_sc_hd__and3_1 c591 (.A(net461),
    .B(net451),
    .C(net462),
    .X(net463));
 sky130_fd_sc_hd__sdfbbn_1 c592 (.CLK_N(clknet_4_6_0_clk),
    .D(net463),
    .RESET_B(net462),
    .SCD(net793),
    .SCE(net460),
    .SET_B(net660),
    .Q(net464));
 sky130_fd_sc_hd__and2_0 c593 (.A(net464),
    .B(net462),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 c594 (.X(net466));
 sky130_fd_sc_hd__clkbuf_1 c595 (.A(net616),
    .X(net467));
 sky130_fd_sc_hd__and3_1 c596 (.A(net370),
    .B(net460),
    .C(net792),
    .X(net468));
 sky130_fd_sc_hd__and3_2 c597 (.A(net319),
    .B(net351),
    .C(net740),
    .X(net469));
 sky130_fd_sc_hd__and3_1 c598 (.A(net185),
    .B(net437),
    .C(net793),
    .X(net470));
 sky130_fd_sc_hd__and2_1 c599 (.A(net332),
    .B(net776),
    .X(net471));
 sky130_fd_sc_hd__sdfbbn_1 c600 (.CLK_N(clknet_4_12_0_clk),
    .D(net468),
    .RESET_B(net265),
    .SCD(net816),
    .SCE(net793),
    .SET_B(net792),
    .Q(net472));
 sky130_fd_sc_hd__and3_1 c601 (.A(net322),
    .B(net715),
    .C(net471),
    .X(net473));
 sky130_fd_sc_hd__and3_1 c602 (.A(net805),
    .B(net471),
    .C(net371),
    .X(net474));
 sky130_fd_sc_hd__and3_1 c603 (.A(net351),
    .B(net109),
    .C(net469),
    .X(net475));
 sky130_fd_sc_hd__and3_1 c604 (.A(net243),
    .B(net702),
    .C(net471),
    .X(net476));
 sky130_fd_sc_hd__and3_2 c605 (.A(net465),
    .B(net185),
    .C(net740),
    .X(net477));
 sky130_fd_sc_hd__and3_1 c606 (.A(net467),
    .B(net471),
    .C(net319),
    .X(net478));
 sky130_fd_sc_hd__and2_0 c607 (.A(net371),
    .B(net77),
    .X(net479));
 sky130_fd_sc_hd__and3_1 c608 (.A(net252),
    .B(net466),
    .C(net837),
    .X(net480));
 sky130_fd_sc_hd__and2_0 c609 (.A(net475),
    .B(net469),
    .X(net481));
 sky130_fd_sc_hd__and3_1 c610 (.A(net236),
    .B(net471),
    .C(net469),
    .X(net482));
 sky130_fd_sc_hd__and3_1 c611 (.A(net715),
    .B(net482),
    .C(net435),
    .X(net483));
 sky130_fd_sc_hd__or4bb_1 c612 (.A(net265),
    .B(net481),
    .C_N(net792),
    .D_N(net477),
    .X(net484));
 sky130_fd_sc_hd__a2111o_1 c613 (.A1(net708),
    .A2(net482),
    .B1(net792),
    .C1(net793),
    .D1(net477),
    .X(net485));
 sky130_fd_sc_hd__sdfbbp_1 c614 (.CLK(clknet_4_3_0_clk),
    .D(net476),
    .RESET_B(net470),
    .SCD(net322),
    .SCE(net484),
    .SET_B(net302),
    .Q(net486));
 sky130_fd_sc_hd__sdfbbn_1 c615 (.CLK_N(clknet_4_12_0_clk),
    .D(net256),
    .RESET_B(net474),
    .SCD(net481),
    .SCE(net261),
    .SET_B(net362),
    .Q(net487));
 sky130_fd_sc_hd__sdfsbp_1 c616 (.CLK(clknet_4_14_0_clk),
    .D(net340),
    .SCD(net384),
    .SCE(net345),
    .SET_B(net867),
    .Q(net738),
    .Q_N(net488));
 sky130_fd_sc_hd__sdfstp_1 c617 (.CLK(clknet_4_14_0_clk),
    .D(net221),
    .SCD(net385),
    .SCE(net735),
    .SET_B(net833),
    .Q(net489));
 sky130_fd_sc_hd__clkbuf_1 c618 (.A(net672),
    .X(net490));
 sky130_fd_sc_hd__sdfstp_1 c619 (.CLK(clknet_4_9_0_clk),
    .D(net457),
    .SCD(net776),
    .SCE(net390),
    .SET_B(net743),
    .Q(net491));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net722),
    .A1(net724),
    .A2(net706),
    .A3(net731),
    .S0(net727),
    .S1(net719),
    .X(net0));
 sky130_fd_sc_hd__and3_1 c620 (.A(net2),
    .B(net45),
    .C(net271),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 c621 (.A(net672),
    .X(net493));
 sky130_fd_sc_hd__sdfxtp_1 c622 (.CLK(clknet_4_13_0_clk),
    .D(net473),
    .SCD(net346),
    .SCE(net302),
    .Q(net494));
 sky130_fd_sc_hd__and3_1 c623 (.A(net384),
    .B(net271),
    .C(net702),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c624 (.A(net493),
    .B(net489),
    .C(net488),
    .X(net747));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net495),
    .A1(net789),
    .A2(net790),
    .A3(net791),
    .S0(net437),
    .S1(net795),
    .X(net496));
 sky130_fd_sc_hd__sdfbbn_1 c626 (.CLK_N(clknet_4_12_0_clk),
    .D(net484),
    .RESET_B(net495),
    .SCD(net741),
    .SCE(net437),
    .SET_B(net271),
    .Q(net497));
 sky130_fd_sc_hd__a2111o_1 c627 (.A1(net390),
    .A2(net869),
    .B1(net45),
    .C1(net387),
    .D1(net776),
    .X(net498));
 sky130_fd_sc_hd__or4bb_1 c628 (.A(net496),
    .B(net490),
    .C_N(net362),
    .D_N(net261),
    .X(net499));
 sky130_fd_sc_hd__sdfxtp_1 c629 (.CLK(clknet_4_11_0_clk),
    .D(net498),
    .SCD(net718),
    .SCE(net765),
    .Q(net737));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net712),
    .A1(net716),
    .A2(net700),
    .A3(net727),
    .S0(net0),
    .S1(net721),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net269),
    .A1(net702),
    .A2(net221),
    .A3(net485),
    .S0(net390),
    .S1(net109),
    .X(net500));
 sky130_fd_sc_hd__and3_1 c631 (.A(net492),
    .B(net744),
    .C(net661),
    .X(net501));
 sky130_fd_sc_hd__dfbbn_1 c632 (.CLK_N(clknet_4_15_0_clk),
    .D(net266),
    .RESET_B(net302),
    .SET_B(net795),
    .Q(net502));
 sky130_fd_sc_hd__and3_1 c633 (.A(net437),
    .B(net398),
    .C(net501),
    .X(net503));
 sky130_fd_sc_hd__dfbbn_1 c634 (.CLK_N(clknet_4_12_0_clk),
    .D(net842),
    .RESET_B(net503),
    .SET_B(net340),
    .Q(net504));
 sky130_fd_sc_hd__a2111o_1 c635 (.A1(net846),
    .A2(net504),
    .B1(net378),
    .C1(net437),
    .D1(net473),
    .X(net505));
 sky130_fd_sc_hd__dfbbp_1 c636 (.CLK(clknet_4_15_0_clk),
    .D(net505),
    .RESET_B(net502),
    .SET_B(net836),
    .Q(net506));
 sky130_fd_sc_hd__sdfstp_1 c637 (.CLK(clknet_4_14_0_clk),
    .D(net499),
    .SCD(net506),
    .SCE(net501),
    .SET_B(net302),
    .Q(net507));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net730),
    .A1(net720),
    .A2(net731),
    .A3(net1),
    .S0(net724),
    .S1(net706),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net706),
    .A1(net682),
    .A2(net711),
    .A3(net679),
    .S0(net734),
    .S1(net705),
    .X(net3));
 sky130_fd_sc_hd__and2_1 c66 (.A(net705),
    .B(net677),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 c660 (.A(net635),
    .X(net508));
 sky130_fd_sc_hd__and2_1 c661 (.A(net305),
    .B(net799),
    .X(net509));
 sky130_fd_sc_hd__and2_0 c662 (.A(net180),
    .B(net421),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_1 c663 (.A(net635),
    .X(net511));
 sky130_fd_sc_hd__and2_1 c664 (.A(net67),
    .B(net822),
    .X(net512));
 sky130_fd_sc_hd__and2_1 c665 (.A(net191),
    .B(net509),
    .X(net513));
 sky130_fd_sc_hd__and2_1 c666 (.A(net511),
    .B(net305),
    .X(net514));
 sky130_fd_sc_hd__and2_1 c667 (.A(net510),
    .B(net799),
    .X(net515));
 sky130_fd_sc_hd__and3_1 c668 (.A(net508),
    .B(net513),
    .C(net305),
    .X(net516));
 sky130_fd_sc_hd__and2_2 c669 (.A(net801),
    .B(net514),
    .X(net517));
 sky130_fd_sc_hd__and2_0 c67 (.A(net682),
    .B(net4),
    .X(net5));
 sky130_fd_sc_hd__dfsbp_1 c670 (.CLK(clknet_4_5_0_clk),
    .D(net295),
    .SET_B(net517),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__dfstp_1 c671 (.CLK(clknet_4_5_0_clk),
    .D(net512),
    .SET_B(net514),
    .Q(net520));
 sky130_fd_sc_hd__dfstp_1 c672 (.CLK(clknet_4_5_0_clk),
    .D(net512),
    .SET_B(net513),
    .Q(net521));
 sky130_fd_sc_hd__and2_0 c673 (.A(net399),
    .B(net521),
    .X(net522));
 sky130_fd_sc_hd__sdfxbp_1 c674 (.CLK(clknet_4_5_0_clk),
    .D(net849),
    .SCD(net410),
    .SCE(net871),
    .Q(net523));
 sky130_fd_sc_hd__sdfxbp_1 c675 (.CLK(clknet_4_5_0_clk),
    .D(net841),
    .SCD(net521),
    .SCE(net410),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__and2_1 c676 (.A(net415),
    .B(net517),
    .X(net526));
 sky130_fd_sc_hd__and2_0 c677 (.A(net508),
    .B(net517),
    .X(net527));
 sky130_fd_sc_hd__and3_1 c678 (.A(net513),
    .B(net518),
    .C(net509),
    .X(net528));
 sky130_fd_sc_hd__and2_1 c679 (.A(net528),
    .B(net524),
    .X(net529));
 sky130_fd_sc_hd__and2_1 c68 (.A(net679),
    .B(net702),
    .X(net6));
 sky130_fd_sc_hd__sdfxtp_1 c680 (.CLK(clknet_4_5_0_clk),
    .D(net527),
    .SCD(net521),
    .SCE(net529),
    .Q(net530));
 sky130_fd_sc_hd__and3_1 c681 (.A(net522),
    .B(net530),
    .C(net794),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net628),
    .X(net532));
 sky130_fd_sc_hd__and2_0 c683 (.A(net531),
    .B(net402),
    .X(net533));
 sky130_fd_sc_hd__and2_0 c684 (.A(net523),
    .B(net402),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 c685 (.A(net850),
    .X(net535));
 sky130_fd_sc_hd__and2_0 c686 (.A(net509),
    .B(net440),
    .X(net536));
 sky130_fd_sc_hd__and3_1 c687 (.A(net315),
    .B(net307),
    .C(net402),
    .X(net537));
 sky130_fd_sc_hd__and3_1 c688 (.A(net533),
    .B(net516),
    .C(net440),
    .X(net538));
 sky130_fd_sc_hd__and2_1 c689 (.A(net98),
    .B(net794),
    .X(net539));
 sky130_fd_sc_hd__and2_1 c69 (.A(net696),
    .B(net700),
    .X(net7));
 sky130_fd_sc_hd__sedfxbp_1 c690 (.CLK(clknet_4_7_0_clk),
    .D(net519),
    .DE(net402),
    .SCD(net538),
    .SCE(net539),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__dfstp_1 c691 (.CLK(clknet_4_7_0_clk),
    .D(net515),
    .SET_B(net538),
    .Q(net542));
 sky130_fd_sc_hd__dlrbn_1 c692 (.D(net538),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net851),
    .Q(net543));
 sky130_fd_sc_hd__and2_0 c693 (.A(net525),
    .B(net542),
    .X(net544));
 sky130_fd_sc_hd__dlrbn_1 c694 (.D(net543),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net538),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__and2_0 c695 (.A(net542),
    .B(net708),
    .X(net547));
 sky130_fd_sc_hd__and2_1 c696 (.A(net328),
    .B(net539),
    .X(net548));
 sky130_fd_sc_hd__dlrbp_1 c697 (.D(net214),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net838),
    .Q(net549));
 sky130_fd_sc_hd__sdfxtp_1 c698 (.CLK(clknet_4_6_0_clk),
    .D(net443),
    .SCD(net547),
    .SCE(net851),
    .Q(net550));
 sky130_fd_sc_hd__dlrbp_1 c699 (.D(net441),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net516),
    .Q(net551));
 sky130_fd_sc_hd__and2_1 c70 (.A(net6),
    .B(net718),
    .X(net8));
 sky130_fd_sc_hd__and2_1 c700 (.A(net549),
    .B(net536),
    .X(net552));
 sky130_fd_sc_hd__or4bb_1 c701 (.A(net440),
    .B(net551),
    .C_N(net552),
    .D_N(net77),
    .X(net553));
 sky130_fd_sc_hd__sedfxbp_1 c702 (.CLK(clknet_4_7_0_clk),
    .D(net553),
    .DE(net519),
    .SCD(net538),
    .SCE(net552),
    .Q(net555),
    .Q_N(net554));
 sky130_fd_sc_hd__or4bb_4 c703 (.A(net550),
    .B(net532),
    .C_N(net540),
    .D_N(net552),
    .X(net556));
 sky130_fd_sc_hd__and2_0 c704 (.A(net537),
    .B(net544),
    .X(net557));
 sky130_fd_sc_hd__or4bb_1 c705 (.A(net717),
    .B(net121),
    .C_N(net517),
    .D_N(net539),
    .X(net558));
 sky130_fd_sc_hd__and3_1 c706 (.A(net552),
    .B(net793),
    .C(net644),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net626),
    .X(net560));
 sky130_fd_sc_hd__and3_1 c708 (.A(net112),
    .B(net539),
    .C(net552),
    .X(net561));
 sky130_fd_sc_hd__and2_0 c709 (.A(net121),
    .B(net454),
    .X(net562));
 sky130_fd_sc_hd__and2_1 c71 (.A(net5),
    .B(net6),
    .X(net9));
 sky130_fd_sc_hd__and2_0 c710 (.A(net516),
    .B(net556),
    .X(net563));
 sky130_fd_sc_hd__and2_0 c711 (.A(net561),
    .B(net793),
    .X(net564));
 sky130_fd_sc_hd__and2_0 c712 (.A(net564),
    .B(net517),
    .X(net565));
 sky130_fd_sc_hd__or4bb_4 c713 (.A(net560),
    .B(net544),
    .C_N(net554),
    .D_N(net556),
    .X(net566));
 sky130_fd_sc_hd__or4bb_1 c714 (.A(net550),
    .B(net566),
    .C_N(net552),
    .D_N(net645),
    .X(net567));
 sky130_fd_sc_hd__or4bb_1 c715 (.A(net454),
    .B(net513),
    .C_N(net456),
    .D_N(net559),
    .X(net568));
 sky130_fd_sc_hd__and2_0 c716 (.A(net456),
    .B(net827),
    .X(net569));
 sky130_fd_sc_hd__and3_1 c717 (.A(net568),
    .B(net826),
    .C(net793),
    .X(net570));
 sky130_fd_sc_hd__or4bb_1 c718 (.A(net514),
    .B(net725),
    .C_N(net825),
    .D_N(net435),
    .X(net571));
 sky130_fd_sc_hd__and3_1 c719 (.A(net562),
    .B(net514),
    .C(net561),
    .X(net572));
 sky130_fd_sc_hd__and2_0 c72 (.A(net719),
    .B(net4),
    .X(net10));
 sky130_fd_sc_hd__and2_0 c720 (.A(net565),
    .B(net567),
    .X(net573));
 sky130_fd_sc_hd__buf_1 c721 (.A(net625),
    .X(net574));
 sky130_fd_sc_hd__sdfbbp_1 c722 (.CLK(clknet_4_7_0_clk),
    .D(net570),
    .RESET_B(net535),
    .SCD(net556),
    .SCE(net526),
    .SET_B(net574),
    .Q(net575));
 sky130_fd_sc_hd__or4bb_1 c723 (.A(net795),
    .B(net301),
    .C_N(net556),
    .D_N(net574),
    .X(net576));
 sky130_fd_sc_hd__and3_1 c724 (.A(net558),
    .B(net575),
    .C(net574),
    .X(net577));
 sky130_fd_sc_hd__and3_1 c725 (.A(net569),
    .B(net576),
    .C(net574),
    .X(net578));
 sky130_fd_sc_hd__sedfxtp_1 c726 (.CLK(clknet_4_6_0_clk),
    .D(net578),
    .DE(net541),
    .SCD(net141),
    .SCE(net674),
    .Q(net579));
 sky130_fd_sc_hd__and3_1 c727 (.A(net534),
    .B(net545),
    .C(net540),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 c728 (.A(net673),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 c729 (.A(net848),
    .X(net582));
 sky130_fd_sc_hd__and2_0 c73 (.A(net10),
    .B(net728),
    .X(net11));
 sky130_fd_sc_hd__sdfbbn_1 c730 (.CLK_N(clknet_4_6_0_clk),
    .D(net141),
    .RESET_B(net446),
    .SCD(net555),
    .SCE(net435),
    .SET_B(net837),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__sdfxtp_1 c731 (.CLK(clknet_4_7_0_clk),
    .D(net563),
    .SCD(net582),
    .SCE(net556),
    .Q(net585));
 sky130_fd_sc_hd__and3_1 c732 (.A(net556),
    .B(net585),
    .C(net435),
    .X(net586));
 sky130_fd_sc_hd__and3_1 c733 (.A(net725),
    .B(net486),
    .C(net517),
    .X(net587));
 sky130_fd_sc_hd__dfbbn_1 c734 (.CLK_N(clknet_4_6_0_clk),
    .D(net483),
    .RESET_B(net480),
    .SET_B(net826),
    .Q(net588));
 sky130_fd_sc_hd__and3_1 c735 (.A(net517),
    .B(net587),
    .C(net581),
    .X(net589));
 sky130_fd_sc_hd__and3_1 c736 (.A(net581),
    .B(net585),
    .C(net725),
    .X(net590));
 sky130_fd_sc_hd__dfbbn_1 c737 (.CLK_N(clknet_4_13_0_clk),
    .D(net361),
    .RESET_B(net826),
    .SET_B(net345),
    .Q(net591));
 sky130_fd_sc_hd__or4bb_4 c738 (.A(net579),
    .B(net580),
    .C_N(net584),
    .D_N(net656),
    .X(net592));
 sky130_fd_sc_hd__or4bb_1 c739 (.A(net586),
    .B(net435),
    .C_N(net526),
    .D_N(net587),
    .X(net593));
 sky130_fd_sc_hd__and2_4 c74 (.A(net1),
    .B(net6),
    .X(net12));
 sky130_fd_sc_hd__and3_1 c740 (.A(net588),
    .B(net446),
    .C(net541),
    .X(net594));
 sky130_fd_sc_hd__or4bb_1 c741 (.A(net559),
    .B(net590),
    .C_N(net593),
    .D_N(net583),
    .X(net595));
 sky130_fd_sc_hd__dfbbp_1 c742 (.CLK(clknet_4_13_0_clk),
    .D(net594),
    .RESET_B(net591),
    .SET_B(net141),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net574),
    .A1(net595),
    .A2(net77),
    .A3(net554),
    .S0(net702),
    .S1(net583),
    .X(net597));
 sky130_fd_sc_hd__and3_1 c744 (.A(net469),
    .B(net592),
    .C(net662),
    .X(net598));
 sky130_fd_sc_hd__a2111o_1 c745 (.A1(net592),
    .A2(net596),
    .B1(net556),
    .C1(net559),
    .D1(net704),
    .X(net599));
 sky130_fd_sc_hd__and3_1 c746 (.A(net598),
    .B(net548),
    .C(net579),
    .X(net600));
 sky130_fd_sc_hd__sdfxbp_1 c747 (.CLK(clknet_4_13_0_clk),
    .D(net600),
    .SCD(net589),
    .SCE(net795),
    .Q(net601));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(net599),
    .A1(net601),
    .A2(net362),
    .A3(net300),
    .S0(net477),
    .S1(net657),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net77),
    .A1(net477),
    .A2(net798),
    .A3(net795),
    .S0(net345),
    .S1(net657),
    .X(net603));
 sky130_fd_sc_hd__and2_0 c75 (.A(net11),
    .B(net6),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net45),
    .A1(net345),
    .A2(net507),
    .A3(net387),
    .S0(net798),
    .S1(clknet_1_1__leaf_net663),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net577),
    .A1(net584),
    .A2(net387),
    .A3(net507),
    .S0(net796),
    .S1(net435),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net478),
    .A1(net362),
    .A2(net487),
    .A3(net77),
    .S0(net796),
    .S1(net584),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net378),
    .A1(net435),
    .A2(net555),
    .A3(net477),
    .S0(net797),
    .S1(clknet_1_0__leaf_net664),
    .X(net607));
 sky130_fd_sc_hd__mux4_2 c754 (.A0(net300),
    .A1(net555),
    .A2(net362),
    .A3(net602),
    .S0(clknet_1_0__leaf_net663),
    .S1(net667),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net109),
    .A1(net472),
    .A2(net798),
    .A3(net665),
    .S0(net666),
    .S1(net668),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net798),
    .A1(net477),
    .A2(net77),
    .A3(clknet_1_1__leaf_net664),
    .S0(net669),
    .S1(net670),
    .X(net610));
 sky130_fd_sc_hd__and2_0 c76 (.A(net13),
    .B(net700),
    .X(net14));
 sky130_fd_sc_hd__and2_1 c77 (.A(net14),
    .B(net6),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c78 (.A(net10),
    .B(net734),
    .X(net16));
 sky130_fd_sc_hd__and2_4 c79 (.A(net12),
    .B(net4),
    .X(net17));
 sky130_fd_sc_hd__and2_4 c80 (.A(net17),
    .B(net16),
    .X(net759));
 sky130_fd_sc_hd__and2_4 c81 (.A(net759),
    .B(net14),
    .X(net18));
 sky130_fd_sc_hd__and2_0 c82 (.A(net7),
    .B(net15),
    .X(net19));
 sky130_fd_sc_hd__and3_1 c83 (.A(net18),
    .B(net759),
    .C(net19),
    .X(net20));
 sky130_fd_sc_hd__and2_4 c84 (.A(net18),
    .B(net7),
    .X(net21));
 sky130_fd_sc_hd__and3_1 c85 (.A(net20),
    .B(net19),
    .C(net21),
    .X(net22));
 sky130_fd_sc_hd__and3_1 c86 (.A(net22),
    .B(net723),
    .C(net21),
    .X(net23));
 sky130_fd_sc_hd__a2111o_1 c87 (.A1(net13),
    .A2(net723),
    .B1(net17),
    .C1(net702),
    .D1(net23),
    .X(net24));
 sky130_fd_sc_hd__and2_1 c88 (.A(net17),
    .B(net5),
    .X(net25));
 sky130_fd_sc_hd__and2_0 c89 (.A(net12),
    .B(net6),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c90 (.A(net11),
    .B(net26),
    .X(net27));
 sky130_fd_sc_hd__and2_1 c91 (.A(net677),
    .B(net759),
    .X(net28));
 sky130_fd_sc_hd__and2_1 c92 (.A(net28),
    .B(net9),
    .X(net29));
 sky130_fd_sc_hd__and2_1 c93 (.A(net26),
    .B(net12),
    .X(net30));
 sky130_fd_sc_hd__and2_0 c94 (.A(net29),
    .B(net9),
    .X(net31));
 sky130_fd_sc_hd__and2_1 c95 (.A(net29),
    .B(net28),
    .X(net32));
 sky130_fd_sc_hd__a2111o_1 c96 (.A1(net27),
    .A2(net30),
    .B1(net28),
    .C1(net31),
    .D1(net25),
    .X(net33));
 sky130_fd_sc_hd__and3_1 c97 (.A(net20),
    .B(net728),
    .C(net702),
    .X(net34));
 sky130_fd_sc_hd__and2_1 c98 (.A(net25),
    .B(net704),
    .X(net35));
 sky130_fd_sc_hd__and2_1 c99 (.A(net677),
    .B(net726),
    .X(net36));
 sky130_fd_sc_hd__sedfxtp_1 merge757 (.CLK(clknet_4_1_0_clk),
    .D(net295),
    .DE(net815),
    .SCD(net302),
    .SCE(net301),
    .Q(net611));
 sky130_fd_sc_hd__sdfxbp_1 merge758 (.CLK(clknet_4_2_0_clk),
    .D(net231),
    .SCD(net112),
    .SCE(net97),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__sdfbbn_1 merge759 (.CLK_N(clknet_4_9_0_clk),
    .D(net847),
    .RESET_B(net362),
    .SCD(net159),
    .SCE(net795),
    .SET_B(net374),
    .Q(net615),
    .Q_N(net614));
 sky130_fd_sc_hd__sdfbbp_1 merge760 (.CLK(clknet_4_6_0_clk),
    .D(net792),
    .RESET_B(net141),
    .SCE(net748),
    .SET_B(net715),
    .Q(net466),
    .Q_N(net616));
 sky130_fd_sc_hd__sedfxtp_1 merge761 (.CLK(clknet_4_2_0_clk),
    .D(net334),
    .DE(net335),
    .SCD(net333),
    .SCE(net337),
    .Q(net618));
 sky130_fd_sc_hd__sdfxtp_1 merge762 (.CLK(clknet_4_0_0_clk),
    .D(net81),
    .SCD(net325),
    .SCE(net861),
    .Q(net619));
 sky130_fd_sc_hd__sdfrbp_1 merge763 (.CLK(clknet_4_9_0_clk),
    .D(net15),
    .RESET_B(net741),
    .SCD(net816),
    .SCE(net756),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__sdfrbp_1 merge764 (.CLK(clknet_4_8_0_clk),
    .D(net146),
    .RESET_B(net804),
    .SCD(net713),
    .SCE(net132),
    .Q(net623),
    .Q_N(net622));
 sky130_fd_sc_hd__sdfrtn_1 merge765 (.CLK_N(clknet_4_9_0_clk),
    .D(net739),
    .RESET_B(net704),
    .SCD(net247),
    .SCE(net124),
    .Q(net624));
 sky130_fd_sc_hd__sdfbbn_1 merge766 (.CLK_N(clknet_4_7_0_clk),
    .D(net346),
    .RESET_B(net571),
    .SCD(net573),
    .SCE(net824),
    .SET_B(net644),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__sdfrtp_1 merge767 (.CLK(clknet_4_10_0_clk),
    .D(net169),
    .RESET_B(net754),
    .SCD(net171),
    .SCE(net708),
    .Q(net627));
 sky130_fd_sc_hd__sdfrtp_1 merge768 (.CLK(clknet_4_5_0_clk),
    .D(net402),
    .RESET_B(net214),
    .SCD(net521),
    .SCE(net529),
    .Q(net628));
 sky130_fd_sc_hd__sdfxtp_1 merge769 (.CLK(clknet_4_11_0_clk),
    .D(net160),
    .SCD(net743),
    .SCE(net271),
    .Q(net629));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net207),
    .A1(net205),
    .A2(net820),
    .A3(net217),
    .S0(net214),
    .S1(net201),
    .X(net630));
 sky130_fd_sc_hd__sdfrtp_1 merge771 (.CLK(clknet_4_6_0_clk),
    .D(net844),
    .RESET_B(net831),
    .SCD(net451),
    .SCE(net354),
    .Q(net631));
 sky130_fd_sc_hd__sdfsbp_1 merge772 (.CLK(clknet_4_1_0_clk),
    .D(net304),
    .SCD(net77),
    .SCE(net195),
    .SET_B(net403),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net447),
    .A1(net485),
    .A2(net718),
    .A3(net354),
    .S0(net479),
    .S1(net776),
    .X(net634));
 sky130_fd_sc_hd__dlrtn_1 merge774 (.D(net420),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net410),
    .Q(net635));
 sky130_fd_sc_hd__sdfsbp_1 merge775 (.CLK(clknet_4_4_0_clk),
    .D(net323),
    .SCD(net321),
    .SCE(net423),
    .SET_B(net792),
    .Q(net637),
    .Q_N(net636));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net557),
    .A1(net526),
    .A2(net469),
    .A3(net572),
    .S0(net346),
    .S1(net556),
    .X(net638));
 sky130_fd_sc_hd__sdfbbn_1 merge777 (.CLK_N(clknet_4_1_0_clk),
    .D(net343),
    .RESET_B(net853),
    .SCD(net304),
    .SCE(net300),
    .SET_B(net67),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__sdfstp_1 merge778 (.CLK(clknet_4_10_0_clk),
    .D(net856),
    .SCD(net221),
    .SCE(net176),
    .SET_B(net140),
    .Q(net641));
 sky130_fd_sc_hd__sdfbbp_1 merge779 (.CLK(clknet_4_2_0_clk),
    .D(net455),
    .RESET_B(net293),
    .SCD(net335),
    .SCE(net237),
    .SET_B(net648),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__dfxbp_1 s780 (.CLK(clknet_4_10_0_clk),
    .D(net179),
    .Q(net779));
 sky130_fd_sc_hd__dfxbp_1 s781 (.CLK(clknet_4_6_0_clk),
    .D(net244),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__dfxtp_1 s782 (.CLK(clknet_4_8_0_clk),
    .D(net263),
    .Q(net646));
 sky130_fd_sc_hd__dfxtp_1 s783 (.CLK(clknet_4_11_0_clk),
    .D(net280),
    .Q(net647));
 sky130_fd_sc_hd__dfxtp_1 s784 (.CLK(clknet_4_11_0_clk),
    .D(net285),
    .Q(net745));
 sky130_fd_sc_hd__dlclkp_1 s785 (.CLK(clknet_4_10_0_clk),
    .GATE(net286),
    .GCLK(net750));
 sky130_fd_sc_hd__dlclkp_2 s786 (.CLK(clknet_4_11_0_clk),
    .GATE(net287),
    .GCLK(net764));
 sky130_fd_sc_hd__dlclkp_4 s787 (.CLK(clknet_4_2_0_clk),
    .GATE(net326),
    .GCLK(net648));
 sky130_fd_sc_hd__dlxbn_1 s788 (.D(net330),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net649));
 sky130_fd_sc_hd__dlxbn_1 s789 (.D(net355),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dlxbp_1 s790 (.D(net356),
    .GATE(clknet_4_3_0_clk),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__dlxtn_1 s791 (.D(net357),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net654));
 sky130_fd_sc_hd__dlxtn_1 s792 (.D(net372),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net655));
 sky130_fd_sc_hd__dlxtn_1 s793 (.D(net377),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net656));
 sky130_fd_sc_hd__dlxtp_1 s794 (.D(net393),
    .GATE(clknet_4_14_0_clk),
    .Q(net657));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s795 (.D(net396),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__dfxbp_1 s796 (.CLK(clknet_4_5_0_clk),
    .D(net439),
    .Q(net658));
 sky130_fd_sc_hd__dfxbp_1 s797 (.CLK(clknet_4_4_0_clk),
    .D(net442),
    .Q(net659));
 sky130_fd_sc_hd__dfxtp_1 s798 (.CLK(clknet_4_6_0_clk),
    .D(net458),
    .Q(net660));
 sky130_fd_sc_hd__dfxtp_1 s799 (.CLK(clknet_4_14_0_clk),
    .D(net500),
    .Q(net661));
 sky130_fd_sc_hd__dfxtp_1 s800 (.CLK(clknet_4_13_0_clk),
    .D(net597),
    .Q(net662));
 sky130_fd_sc_hd__dlclkp_1 s801 (.CLK(clknet_4_15_0_clk),
    .GATE(net603),
    .GCLK(net663));
 sky130_fd_sc_hd__dlclkp_2 s802 (.CLK(clknet_4_15_0_clk),
    .GATE(net604),
    .GCLK(net664));
 sky130_fd_sc_hd__dlclkp_4 s803 (.CLK(clknet_4_15_0_clk),
    .GATE(net605),
    .GCLK(net665));
 sky130_fd_sc_hd__dlxbn_1 s804 (.D(net606),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__dlxbn_1 s805 (.D(net607),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net667));
 sky130_fd_sc_hd__dlxbp_1 s806 (.D(net608),
    .GATE(clknet_4_15_0_clk),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__dlxtn_1 s807 (.D(net609),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net670));
 sky130_fd_sc_hd__dlxtn_2 s808 (.D(net610),
    .GATE_N(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlxtn_1 s809 (.D(net630),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net671));
 sky130_fd_sc_hd__dlxtp_1 s810 (.D(net634),
    .GATE(clknet_4_13_0_clk),
    .Q(net672));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s811 (.D(net638),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net673));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net675));
 sky130_fd_sc_hd__buf_1 input4 (.A(in11),
    .X(net676));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net677));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net679));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net680));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net681));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(in17),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net683));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net684));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(in2),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in20),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in22),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in26),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net695));
 sky130_fd_sc_hd__buf_1 input24 (.A(in3),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in32),
    .X(net699));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net701));
 sky130_fd_sc_hd__buf_4 input30 (.A(in35),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net703));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net704));
 sky130_fd_sc_hd__buf_2 input33 (.A(in38),
    .X(net705));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in4),
    .X(net707));
 sky130_fd_sc_hd__buf_4 input36 (.A(in40),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net710));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in44),
    .X(net712));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net714));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net715));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net716));
 sky130_fd_sc_hd__buf_2 input45 (.A(in49),
    .X(net717));
 sky130_fd_sc_hd__buf_4 input46 (.A(in5),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(in50),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(in51),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(in52),
    .X(net721));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net722));
 sky130_fd_sc_hd__buf_1 input51 (.A(in54),
    .X(net723));
 sky130_fd_sc_hd__buf_6 input52 (.A(in55),
    .X(net724));
 sky130_fd_sc_hd__buf_2 input53 (.A(in56),
    .X(net725));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net726));
 sky130_fd_sc_hd__buf_8 input55 (.A(in58),
    .X(net727));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net728));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net729));
 sky130_fd_sc_hd__buf_1 input58 (.A(in60),
    .X(net730));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(in7),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in8),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(in9),
    .X(net734));
 sky130_fd_sc_hd__buf_2 output63 (.A(net735),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net736),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net737),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net738),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net739),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net740),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net741),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net742),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net743),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output72 (.A(net744),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net745),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net746),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net747),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net748),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net749),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net750),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output79 (.A(net751),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output80 (.A(net752),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output81 (.A(net753),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output82 (.A(net754),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output83 (.A(net755),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output84 (.A(net756),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net757),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output86 (.A(net758),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output87 (.A(net759),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output88 (.A(net760),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output89 (.A(net761),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output90 (.A(net762),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output91 (.A(net763),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(clknet_1_1__leaf_net764),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output93 (.A(net765),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output94 (.A(net766),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output95 (.A(net767),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output96 (.A(net768),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output97 (.A(net769),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output98 (.A(net770),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output99 (.A(net771),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output100 (.A(net794),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output101 (.A(net773),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net774),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output103 (.A(net775),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output104 (.A(net776),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output105 (.A(net777),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output106 (.A(net778),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output107 (.A(net779),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output108 (.A(net780),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output109 (.A(net781),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output110 (.A(net782),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output111 (.A(net783),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output112 (.A(net784),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output113 (.A(net785),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output114 (.A(net786),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net787),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output116 (.A(net788),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output117 (.A(net789),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output118 (.A(net790),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output119 (.A(net791),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net327),
    .X(net792));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net446),
    .X(net793));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net772),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net772),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net664 (.A(net664),
    .X(clknet_0_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_0__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net664 (.A(clknet_0_net664),
    .X(clknet_1_1__leaf_net664));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net663 (.A(net663),
    .X(clknet_0_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_0__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net663 (.A(clknet_0_net663),
    .X(clknet_1_1__leaf_net663));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net764 (.A(net764),
    .X(clknet_0_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_0__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net764 (.A(clknet_0_net764),
    .X(clknet_1_1__leaf_net764));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net750 (.A(net750),
    .X(clknet_0_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_0__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_1__leaf_net750));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net602),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net602),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net602),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net83),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net799),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net799),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net24),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net23),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net22),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net813),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net73),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net293),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net293),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net816),
    .X(net817));
 sky130_fd_sc_hd__buf_2 rebuffer23 (.A(net817),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net159),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net200),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net820),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net200),
    .X(net822));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer28 (.A(net200),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer29 (.A(net566),
    .X(net824));
 sky130_fd_sc_hd__bufbuf_8 rebuffer30 (.A(net824),
    .X(net825));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer31 (.A(net825),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net826),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net759),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net75),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net646),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net345),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net632),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net383),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net275),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net359),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net657),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net656),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net546),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net348),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net368),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net422),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net497),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net238),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net430),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net382),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net494),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net149),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net673),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net520),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net628),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net542),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net161),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net349),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net262),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net148),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net274),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net251),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net328),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net659),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net647),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net311),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net620),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net164),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net416),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net379),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net232),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net776),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net235),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net491),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net652),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net518),
    .X(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_D_N (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_D1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge758_SCD (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_D_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_D1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_RESET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_D (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_C (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_SCD (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCE (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SET_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCE (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_RESET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_D (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_SCD (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_SCD (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCD (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCE (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Q (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCD (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_D (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_D_N (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_D_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SCE (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_Q_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_D (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_C (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCE (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_C (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_C (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_SCD (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_RESET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCE (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_S1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_SCE (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_SET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCE (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SCD (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_RESET_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_C (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_SCD (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_D1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_RESET_B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SET_B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCD (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCE (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SET_B (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_S0 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_D (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCE (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCD (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_SCE (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_RESET_B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_C_N (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SET_B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_C (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SET_B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_B1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_C1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_C (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_Q (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_SCE (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_D_N (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_X (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_C1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SCE (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_C (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_C (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_X (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_D1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_D_N (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_SET_B (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_X (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_SET_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_C (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C_N (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_SET_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_SCD (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_Q (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_Q_N (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_D1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_Q (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D_N (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_s794_Q (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_C (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_SCD (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_D_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_RESET_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_SCE (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge758_SCE (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCE (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_C (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_SCD (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_C (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_C1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_C (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_RESET_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_D1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_D (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCE (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_C (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_SET_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCD (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_C (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_RESET_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_SCE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S0 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_D1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_C (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_RESET_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SCE (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_D (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_C (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_C (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_X (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_RESET_B (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SCD (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_SCD (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_Q (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_SCD (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SET_B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_SCE (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCD (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCE (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_RESET_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_SCD (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_SCE (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_C_N (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SCD (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_X (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCE (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_RESET_B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCE (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_RESET_B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCE (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_D1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SCD (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCE (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_D1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SCE (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SET_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_C (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SCE (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge760_D (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_B1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SET_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_C (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_SET_B (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_SCE (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_SCE (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_C (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_C (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_C1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_C (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_C (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_SCD (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C_N (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_C (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_C (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_D_N (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_SCE (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCE (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_SET_B (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_D1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s788_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s797_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_D (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_SCE (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold59_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SET_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net84),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net872),
    .X(net873));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer37 (.A(net873),
    .X(net874));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer38 (.A(net872),
    .X(net875));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
