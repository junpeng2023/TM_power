module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net632;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net782;
 wire clknet_1_0__leaf_net782;
 wire clknet_1_1__leaf_net782;
 wire clknet_0_net449;
 wire clknet_1_0__leaf_net449;
 wire clknet_1_1__leaf_net449;
 wire clknet_0_net243;
 wire clknet_1_0__leaf_net243;
 wire clknet_1_1__leaf_net243;
 wire clknet_0_net257;
 wire clknet_1_0__leaf_net257;
 wire clknet_1_1__leaf_net257;
 wire clknet_0_net262;
 wire clknet_1_0__leaf_net262;
 wire clknet_1_1__leaf_net262;
 wire clknet_0_net269;
 wire clknet_1_0__leaf_net269;
 wire clknet_1_1__leaf_net269;
 wire clknet_0_net854;
 wire clknet_1_0__leaf_net854;
 wire clknet_1_1__leaf_net854;
 wire clknet_0_net894;
 wire clknet_1_0__leaf_net894;
 wire clknet_1_1__leaf_net894;
 wire clknet_0_net874;
 wire clknet_1_0__leaf_net874;
 wire clknet_1_1__leaf_net874;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net265;
 wire clknet_1_0__leaf_net265;
 wire clknet_1_1__leaf_net265;
 wire clknet_0_net781;
 wire clknet_1_0__leaf_net781;
 wire clknet_1_1__leaf_net781;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire clknet_0_net423;
 wire clknet_1_0__leaf_net423;
 wire clknet_1_1__leaf_net423;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net537;
 wire clknet_1_0__leaf_net537;
 wire clknet_1_1__leaf_net537;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net548;
 wire clknet_1_0__leaf_net548;
 wire clknet_1_1__leaf_net548;
 wire clknet_0_net538;
 wire clknet_1_0__leaf_net538;
 wire clknet_1_1__leaf_net538;
 wire clknet_0_net762;
 wire clknet_1_0__leaf_net762;
 wire clknet_1_1__leaf_net762;
 wire clknet_0_net433;
 wire clknet_1_0__leaf_net433;
 wire clknet_1_1__leaf_net433;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net474;
 wire clknet_1_0__leaf_net474;
 wire clknet_1_1__leaf_net474;
 wire clknet_0_net761;
 wire clknet_1_0__leaf_net761;
 wire clknet_1_1__leaf_net761;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net428;
 wire clknet_1_0__leaf_net428;
 wire clknet_1_1__leaf_net428;
 wire clknet_0_net780;
 wire clknet_1_0__leaf_net780;
 wire clknet_1_1__leaf_net780;
 wire clknet_0_net431;
 wire clknet_1_0__leaf_net431;
 wire clknet_1_1__leaf_net431;
 wire clknet_0_net425;
 wire clknet_1_0__leaf_net425;
 wire clknet_1_1__leaf_net425;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net760;
 wire clknet_1_0__leaf_net760;
 wire clknet_1_1__leaf_net760;
 wire clknet_0_net550;
 wire clknet_1_0__leaf_net550;
 wire clknet_1_1__leaf_net550;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net545;
 wire clknet_1_0__leaf_net545;
 wire clknet_1_1__leaf_net545;
 wire clknet_0_net551;
 wire clknet_1_0__leaf_net551;
 wire clknet_1_1__leaf_net551;
 wire clknet_0_net741;
 wire clknet_1_0__leaf_net741;
 wire clknet_1_1__leaf_net741;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net724;
 wire clknet_1_0__leaf_net724;
 wire clknet_1_1__leaf_net724;
 wire clknet_0_net521;
 wire clknet_1_0__leaf_net521;
 wire clknet_1_1__leaf_net521;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net520;
 wire clknet_1_0__leaf_net520;
 wire clknet_1_1__leaf_net520;
 wire clknet_0_net528;
 wire clknet_1_0__leaf_net528;
 wire clknet_1_1__leaf_net528;
 wire clknet_0_net518;
 wire clknet_1_0__leaf_net518;
 wire clknet_1_1__leaf_net518;
 wire clknet_0_net513;
 wire clknet_1_0__leaf_net513;
 wire clknet_1_1__leaf_net513;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net529;
 wire clknet_1_0__leaf_net529;
 wire clknet_1_1__leaf_net529;
 wire clknet_0_net535;
 wire clknet_1_0__leaf_net535;
 wire clknet_1_1__leaf_net535;
 wire clknet_0_net591;
 wire clknet_1_0__leaf_net591;
 wire clknet_1_1__leaf_net591;
 wire clknet_0_net531;
 wire clknet_1_0__leaf_net531;
 wire clknet_1_1__leaf_net531;
 wire clknet_0_net519;
 wire clknet_1_0__leaf_net519;
 wire clknet_1_1__leaf_net519;
 wire clknet_0_net408;
 wire clknet_1_0__leaf_net408;
 wire clknet_1_1__leaf_net408;
 wire clknet_0_net526;
 wire clknet_1_0__leaf_net526;
 wire clknet_1_1__leaf_net526;
 wire clknet_0_net406;
 wire clknet_1_0__leaf_net406;
 wire clknet_1_1__leaf_net406;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net486;
 wire clknet_1_0__leaf_net486;
 wire clknet_1_1__leaf_net486;
 wire clknet_0_net620;
 wire clknet_1_0__leaf_net620;
 wire clknet_1_1__leaf_net620;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net416;
 wire clknet_1_0__leaf_net416;
 wire clknet_1_1__leaf_net416;
 wire clknet_0_net394;
 wire clknet_1_0__leaf_net394;
 wire clknet_1_1__leaf_net394;
 wire clknet_0_net706;
 wire clknet_1_0__leaf_net706;
 wire clknet_1_1__leaf_net706;
 wire clknet_0_net419;
 wire clknet_1_0__leaf_net419;
 wire clknet_1_1__leaf_net419;
 wire clknet_0_net692;
 wire clknet_1_0__leaf_net692;
 wire clknet_1_1__leaf_net692;
 wire clknet_0_net361;
 wire clknet_1_0__leaf_net361;
 wire clknet_1_1__leaf_net361;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net362;
 wire clknet_1_0__leaf_net362;
 wire clknet_1_1__leaf_net362;
 wire clknet_0_net371;
 wire clknet_1_0__leaf_net371;
 wire clknet_1_1__leaf_net371;
 wire clknet_0_net860;
 wire clknet_1_0__leaf_net860;
 wire clknet_1_1__leaf_net860;
 wire clknet_0_net862;
 wire clknet_1_0__leaf_net862;
 wire clknet_1_1__leaf_net862;
 wire clknet_0_net377;
 wire clknet_1_0__leaf_net377;
 wire clknet_1_1__leaf_net377;
 wire clknet_0_net861;
 wire clknet_1_0__leaf_net861;
 wire clknet_1_1__leaf_net861;
 wire clknet_0_net364;
 wire clknet_1_0__leaf_net364;
 wire clknet_1_1__leaf_net364;
 wire clknet_0_net873;
 wire clknet_1_0__leaf_net873;
 wire clknet_1_1__leaf_net873;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net899;
 wire clknet_1_0__leaf_net899;
 wire clknet_1_1__leaf_net899;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net171;
 wire clknet_1_0__leaf_net171;
 wire clknet_1_1__leaf_net171;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;

 sky130_fd_sc_hd__a21bo_1 c100 (.A1(net3),
    .A2(net22),
    .B1_N(net28),
    .X(net37));
 sky130_fd_sc_hd__a31o_4 c101 (.A1(net26),
    .A2(net36),
    .A3(net28),
    .B1(net930),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net31),
    .A1(net6),
    .A2(net29),
    .A3(net38),
    .S0(net805),
    .S1(net28),
    .X(net887));
 sky130_fd_sc_hd__a21bo_1 c103 (.A1(net36),
    .A2(net29),
    .B1_N(net38),
    .X(net39));
 sky130_fd_sc_hd__a21bo_2 c104 (.A1(net39),
    .A2(net35),
    .B1_N(net37),
    .X(net40));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net7),
    .A2(net30),
    .B1_N(net31),
    .X(net41));
 sky130_fd_sc_hd__a21bo_1 c106 (.A1(net33),
    .A2(net41),
    .B1_N(net38),
    .X(net42));
 sky130_fd_sc_hd__a21bo_1 c107 (.A1(net16),
    .A2(net805),
    .B1_N(net41),
    .X(net43));
 sky130_fd_sc_hd__a21bo_1 c108 (.A1(net42),
    .A2(net43),
    .B1_N(net32),
    .X(net44));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net43),
    .A1(net41),
    .A2(net887),
    .A3(net44),
    .S0(net845),
    .S1(net25),
    .X(net881));
 sky130_fd_sc_hd__xnor2_4 c110 (.A(net36),
    .B(net938),
    .Y(net893));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net792),
    .B(net945),
    .Y(net890));
 sky130_fd_sc_hd__xnor2_4 c112 (.A(net930),
    .B(net938),
    .Y(net45));
 sky130_fd_sc_hd__xnor2_4 c113 (.A(net943),
    .B(net893),
    .Y(net46));
 sky130_fd_sc_hd__a21bo_1 c114 (.A1(net893),
    .A2(net943),
    .B1_N(net43),
    .X(net47));
 sky130_fd_sc_hd__xnor2_4 c115 (.A(net828),
    .B(net46),
    .Y(net48));
 sky130_fd_sc_hd__xnor2_4 c116 (.A(net40),
    .B(net25),
    .Y(net49));
 sky130_fd_sc_hd__xnor2_2 c117 (.A(net0),
    .B(net49),
    .Y(net868));
 sky130_fd_sc_hd__a41o_1 c118 (.A1(net47),
    .A2(net944),
    .A3(net839),
    .A4(net868),
    .B1(net40),
    .X(net888));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net46),
    .B(net922),
    .Y(net50));
 sky130_fd_sc_hd__xnor2_4 c120 (.A(net45),
    .B(net49),
    .Y(net51));
 sky130_fd_sc_hd__xnor2_1 c121 (.A(net43),
    .B(net45),
    .Y(net878));
 sky130_fd_sc_hd__xnor2_4 c122 (.A(net48),
    .B(net51),
    .Y(net871));
 sky130_fd_sc_hd__a31o_1 c123 (.A1(net33),
    .A2(net890),
    .A3(net46),
    .B1(net25),
    .X(net52));
 sky130_fd_sc_hd__a41o_2 c124 (.A1(net52),
    .A2(net871),
    .A3(net48),
    .A4(net50),
    .B1(net939),
    .X(net896));
 sky130_fd_sc_hd__a21bo_1 c125 (.A1(net51),
    .A2(net937),
    .B1_N(net896),
    .X(net53));
 sky130_fd_sc_hd__a41o_1 c126 (.A1(net35),
    .A2(net871),
    .A3(net896),
    .A4(net52),
    .B1(net888),
    .X(net54));
 sky130_fd_sc_hd__a41o_1 c127 (.A1(net50),
    .A2(net878),
    .A3(net52),
    .A4(net896),
    .B1(net54),
    .X(net55));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net834),
    .A2(net52),
    .A3(net55),
    .A4(net871),
    .B1(net47),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net53),
    .A1(net52),
    .A2(net940),
    .A3(net50),
    .S0(net896),
    .S1(net55),
    .X(net57));
 sky130_fd_sc_hd__a41o_1 c130 (.A1(net53),
    .A2(net36),
    .A3(net28),
    .A4(net657),
    .B1(net700),
    .X(net855));
 sky130_fd_sc_hd__a41o_1 c131 (.A1(net55),
    .A2(net871),
    .A3(net855),
    .B1(net700),
    .X(net58));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net800),
    .B(net820),
    .Y(net59));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net788),
    .B(net793),
    .Y(net60));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net59),
    .B(net790),
    .Y(net61));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net632),
    .B(net796),
    .Y(net62));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net62),
    .B(net793),
    .Y(net63));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net61),
    .B(net790),
    .Y(net64));
 sky130_fd_sc_hd__a31o_4 c138 (.A1(net63),
    .A2(net62),
    .A3(net800),
    .B1(net809),
    .X(net65));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net60),
    .B(net799),
    .Y(net66));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net65),
    .B(net809),
    .Y(net67));
 sky130_fd_sc_hd__a31o_1 c141 (.A1(net63),
    .A2(net64),
    .A3(net66),
    .B1(net65),
    .X(net68));
 sky130_fd_sc_hd__xnor2_4 c142 (.A(net67),
    .B(net787),
    .Y(net69));
 sky130_fd_sc_hd__a21bo_1 c143 (.A1(net68),
    .A2(net64),
    .B1_N(net69),
    .X(net70));
 sky130_fd_sc_hd__a41o_2 c144 (.A1(net65),
    .A2(net792),
    .A3(net70),
    .A4(net66),
    .B1(net68),
    .X(net71));
 sky130_fd_sc_hd__a41o_2 c145 (.A1(net70),
    .A2(net820),
    .A3(net61),
    .A4(net71),
    .B1(net59),
    .X(net72));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net790),
    .A2(net66),
    .A3(net793),
    .A4(net789),
    .B1(net820),
    .X(net73));
 sky130_fd_sc_hd__a41o_4 c147 (.A1(net72),
    .A2(net73),
    .A3(net67),
    .A4(net64),
    .B1(net71),
    .X(net74));
 sky130_fd_sc_hd__a21bo_1 c148 (.A1(net820),
    .A2(net65),
    .B1_N(net67),
    .X(net75));
 sky130_fd_sc_hd__a41o_2 c149 (.A1(net70),
    .A2(net74),
    .A3(net60),
    .A4(net67),
    .B1(net929),
    .X(net76));
 sky130_fd_sc_hd__a41o_4 c150 (.A1(net795),
    .A2(net69),
    .A3(net929),
    .A4(net76),
    .B1(net66),
    .X(net77));
 sky130_fd_sc_hd__a21bo_4 c151 (.A1(net929),
    .A2(net76),
    .B1_N(net799),
    .X(net78));
 sky130_fd_sc_hd__a41o_4 c152 (.A1(net74),
    .A2(net69),
    .A3(net62),
    .A4(net73),
    .B1(net75),
    .X(net79));
 sky130_fd_sc_hd__a41o_4 c153 (.A1(net792),
    .A2(net78),
    .A3(net77),
    .A4(net76),
    .B1(net65),
    .X(net80));
 sky130_fd_sc_hd__xnor2_1 c154 (.A(net71),
    .B(net805),
    .Y(net81));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net803),
    .B(net74),
    .Y(net82));
 sky130_fd_sc_hd__a31o_2 c156 (.A1(net802),
    .A2(net82),
    .A3(net817),
    .B1(net815),
    .X(net83));
 sky130_fd_sc_hd__xnor2_1 c157 (.A(net822),
    .B(net82),
    .Y(net84));
 sky130_fd_sc_hd__a21bo_1 c158 (.A1(net83),
    .A2(net78),
    .B1_N(net82),
    .X(net85));
 sky130_fd_sc_hd__a21bo_1 c159 (.A1(net810),
    .A2(net804),
    .B1_N(net916),
    .X(net86));
 sky130_fd_sc_hd__a31o_4 c160 (.A1(net59),
    .A2(net61),
    .A3(net916),
    .B1(net82),
    .X(net87));
 sky130_fd_sc_hd__xnor2_1 c161 (.A(net82),
    .B(net71),
    .Y(net88));
 sky130_fd_sc_hd__mux4_2 c162 (.A0(net818),
    .A1(net72),
    .A2(net83),
    .A3(net87),
    .S0(net60),
    .S1(net916),
    .X(net89));
 sky130_fd_sc_hd__a21bo_4 c163 (.A1(net89),
    .A2(net812),
    .B1_N(net916),
    .X(net90));
 sky130_fd_sc_hd__a21bo_1 c164 (.A1(net88),
    .A2(net831),
    .B1_N(net72),
    .X(net91));
 sky130_fd_sc_hd__a21bo_1 c165 (.A1(net91),
    .A2(net794),
    .B1_N(net87),
    .X(net92));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net815),
    .A1(net71),
    .A2(net808),
    .A3(net797),
    .S0(net79),
    .S1(net917),
    .X(net93));
 sky130_fd_sc_hd__a21bo_1 c167 (.A1(net93),
    .A2(net83),
    .B1_N(net917),
    .X(net94));
 sky130_fd_sc_hd__a41o_2 c168 (.A1(net92),
    .A2(net93),
    .A3(net90),
    .A4(net805),
    .B1(net916),
    .X(net95));
 sky130_fd_sc_hd__a21bo_1 c169 (.A1(net82),
    .A2(net95),
    .B1_N(net916),
    .X(net96));
 sky130_fd_sc_hd__a31o_4 c170 (.A1(net96),
    .A2(net94),
    .A3(net95),
    .B1(net64),
    .X(net97));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net95),
    .A1(net97),
    .A2(net82),
    .A3(net86),
    .S0(net93),
    .S1(net96),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net816),
    .A1(net94),
    .A2(net808),
    .A3(net98),
    .S0(net95),
    .S1(net89),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net81),
    .A1(net93),
    .A2(net98),
    .A3(net86),
    .S0(net64),
    .S1(net916),
    .X(net100));
 sky130_fd_sc_hd__a21bo_4 c174 (.A1(net819),
    .A2(net95),
    .B1_N(net98),
    .X(net856));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net99),
    .A1(net94),
    .A2(net93),
    .A3(net97),
    .S0(net98),
    .S1(net916),
    .X(net101));
 sky130_fd_sc_hd__xnor2_4 c176 (.A(net80),
    .B(net798),
    .Y(net102));
 sky130_fd_sc_hd__xnor2_4 c177 (.A(net829),
    .B(net832),
    .Y(net103));
 sky130_fd_sc_hd__a31o_1 c178 (.A1(net824),
    .A2(net102),
    .A3(net80),
    .B1(net843),
    .X(net104));
 sky130_fd_sc_hd__xnor2_4 c179 (.A(net87),
    .B(net66),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_4 c180 (.A(net102),
    .B(net105),
    .Y(net106));
 sky130_fd_sc_hd__a31o_2 c181 (.A1(net72),
    .A2(net843),
    .A3(net813),
    .B1(net808),
    .X(net107));
 sky130_fd_sc_hd__a31o_1 c182 (.A1(net69),
    .A2(net837),
    .A3(net87),
    .B1(net107),
    .X(net108));
 sky130_fd_sc_hd__xnor2_4 c183 (.A(net103),
    .B(net824),
    .Y(net109));
 sky130_fd_sc_hd__a31o_4 c184 (.A1(net84),
    .A2(net838),
    .A3(net103),
    .B1(net107),
    .X(net110));
 sky130_fd_sc_hd__a21bo_2 c185 (.A1(net104),
    .A2(net107),
    .B1_N(net60),
    .X(net111));
 sky130_fd_sc_hd__xnor2_4 c186 (.A(net979),
    .B(net111),
    .Y(net112));
 sky130_fd_sc_hd__mux4_2 c187 (.A0(net111),
    .A1(net937),
    .A2(net109),
    .A3(net829),
    .S0(net107),
    .S1(net839),
    .X(net113));
 sky130_fd_sc_hd__xnor2_2 c188 (.A(net60),
    .B(net105),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_1 c189 (.A(net113),
    .B(net979),
    .Y(net115));
 sky130_fd_sc_hd__xnor2_1 c190 (.A(net115),
    .B(net910),
    .Y(net116));
 sky130_fd_sc_hd__clkbuf_1 c191 (.A(net687),
    .X(net117));
 sky130_fd_sc_hd__xnor2_4 c192 (.A(net910),
    .B(net109),
    .Y(net118));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net838),
    .A1(net109),
    .A2(net118),
    .A3(net832),
    .S0(net112),
    .S1(net115),
    .X(net119));
 sky130_fd_sc_hd__a31o_1 c194 (.A1(net118),
    .A2(net111),
    .A3(net116),
    .B1(net117),
    .X(net120));
 sky130_fd_sc_hd__mux4_2 c195 (.A0(net799),
    .A1(net116),
    .A2(net119),
    .A3(net86),
    .S0(net113),
    .S1(net910),
    .X(net121));
 sky130_fd_sc_hd__xnor2_4 c196 (.A(net121),
    .B(net118),
    .Y(net122));
 sky130_fd_sc_hd__a31o_1 c197 (.A1(net117),
    .A2(net109),
    .A3(net122),
    .B1(net87),
    .X(net123));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net806),
    .A2(net856),
    .B1_N(net119),
    .X(net124));
 sky130_fd_sc_hd__buf_1 c199 (.A(net687),
    .X(net125));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net76),
    .A2(net19),
    .B1_N(net90),
    .X(net126));
 sky130_fd_sc_hd__buf_1 c201 (.A(net687),
    .X(net127));
 sky130_fd_sc_hd__a21bo_2 c202 (.A1(net24),
    .A2(net108),
    .B1_N(net126),
    .X(net128));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net125),
    .A2(net114),
    .B1_N(net127),
    .X(net129));
 sky130_fd_sc_hd__a21bo_1 c204 (.A1(net108),
    .A2(net922),
    .B1_N(net106),
    .X(net130));
 sky130_fd_sc_hd__a21bo_2 c205 (.A1(net126),
    .A2(net127),
    .B1_N(net844),
    .X(net131));
 sky130_fd_sc_hd__a21bo_1 c206 (.A1(net15),
    .A2(net129),
    .B1_N(net24),
    .X(net132));
 sky130_fd_sc_hd__a21bo_1 c207 (.A1(net5),
    .A2(net131),
    .B1_N(net64),
    .X(net133));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(net133),
    .A2(net125),
    .B1_N(net127),
    .X(net134));
 sky130_fd_sc_hd__mux4_2 c209 (.A0(net109),
    .A1(net134),
    .A2(net12),
    .A3(net112),
    .S0(net125),
    .S1(net6),
    .X(net135));
 sky130_fd_sc_hd__a31o_1 c210 (.A1(net129),
    .A2(net134),
    .A3(net119),
    .B1(net130),
    .X(net136));
 sky130_fd_sc_hd__a21bo_2 c211 (.A1(net127),
    .A2(net856),
    .B1_N(net12),
    .X(net137));
 sky130_fd_sc_hd__a31o_2 c212 (.A1(net136),
    .A2(net128),
    .A3(net90),
    .B1(net832),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net813),
    .A1(net122),
    .A2(net138),
    .A3(net73),
    .S0(net109),
    .S1(net78),
    .X(net139));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(net114),
    .A2(net905),
    .A3(net23),
    .A4(net137),
    .B1(net701),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net131),
    .A1(net120),
    .A2(net15),
    .A3(net126),
    .S0(net813),
    .S1(net687),
    .X(net141));
 sky130_fd_sc_hd__a31o_1 c216 (.A1(net141),
    .A2(net839),
    .A3(net15),
    .B1(net701),
    .X(net142));
 sky130_fd_sc_hd__a41o_1 c217 (.A1(net12),
    .A2(net134),
    .A3(net90),
    .A4(net125),
    .B1(net701),
    .X(net143));
 sky130_fd_sc_hd__a41o_1 c218 (.A1(net142),
    .A2(net126),
    .A3(net137),
    .A4(net130),
    .B1(net687),
    .X(net144));
 sky130_fd_sc_hd__sdfrbp_2 c219 (.CLK(clknet_4_13_0_clk),
    .D(net143),
    .RESET_B(net137),
    .SCD(net687),
    .SCE(net702),
    .Q(net895),
    .Q_N(net145));
 sky130_fd_sc_hd__xnor2_2 c220 (.A(net9),
    .B(net881),
    .Y(net146));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(net44),
    .B(net844),
    .Y(net147));
 sky130_fd_sc_hd__xnor2_2 c222 (.A(net131),
    .B(net73),
    .Y(net900));
 sky130_fd_sc_hd__xnor2_1 c223 (.A(net847),
    .B(net44),
    .Y(net148));
 sky130_fd_sc_hd__xnor2_1 c224 (.A(net6),
    .B(net980),
    .Y(net149));
 sky130_fd_sc_hd__xnor2_1 c225 (.A(net63),
    .B(net145),
    .Y(net150));
 sky130_fd_sc_hd__xnor2_4 c226 (.A(net79),
    .B(net145),
    .Y(net151));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(net146),
    .A2(net804),
    .B1_N(net151),
    .X(net152));
 sky130_fd_sc_hd__xnor2_1 c228 (.A(net151),
    .B(net134),
    .Y(net153));
 sky130_fd_sc_hd__xnor2_1 c229 (.A(net147),
    .B(net44),
    .Y(net154));
 sky130_fd_sc_hd__xnor2_4 c230 (.A(net980),
    .B(net907),
    .Y(net155));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net844),
    .A2(net151),
    .B1_N(net155),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net155),
    .A1(net131),
    .A2(net112),
    .A3(net907),
    .S0(net151),
    .S1(net906),
    .X(net157));
 sky130_fd_sc_hd__mux4_2 c233 (.A0(net156),
    .A1(net906),
    .A2(net147),
    .A3(net28),
    .S0(net37),
    .S1(net907),
    .X(net158));
 sky130_fd_sc_hd__a21bo_4 c234 (.A1(net37),
    .A2(net151),
    .B1_N(net155),
    .X(net159));
 sky130_fd_sc_hd__a21bo_1 c235 (.A1(net789),
    .A2(net156),
    .B1_N(net155),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net90),
    .A1(net844),
    .A2(net904),
    .A3(net156),
    .S0(net151),
    .S1(net146),
    .X(net161));
 sky130_fd_sc_hd__a21bo_1 c237 (.A1(net155),
    .A2(net151),
    .B1_N(net904),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 c238 (.A(net950),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net160),
    .A1(net153),
    .A2(net158),
    .A3(net162),
    .S0(net156),
    .S1(net941),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 c240 (.A(net662),
    .X(net165));
 sky130_fd_sc_hd__a41o_1 c241 (.A1(net165),
    .A2(net905),
    .A3(net156),
    .A4(net955),
    .B1(net662),
    .X(net166));
 sky130_fd_sc_hd__a21bo_1 c242 (.A1(net64),
    .A2(net890),
    .B1_N(net871),
    .X(net875));
 sky130_fd_sc_hd__buf_1 c243 (.A(clknet_1_0__leaf_net898),
    .X(net899));
 sky130_fd_sc_hd__a21bo_1 c244 (.A1(net28),
    .A2(net881),
    .B1_N(net702),
    .X(net167));
 sky130_fd_sc_hd__sdfrbp_1 c245 (.CLK(clknet_4_15_0_clk),
    .D(net132),
    .RESET_B(net893),
    .SCD(net137),
    .SCE(net656),
    .Q(net169),
    .Q_N(net168));
 sky130_fd_sc_hd__a31o_1 c246 (.A1(net128),
    .A2(net922),
    .A3(net657),
    .B1(net897),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c247 (.A(clknet_1_0__leaf_net898),
    .X(net879));
 sky130_fd_sc_hd__a21bo_1 c248 (.A1(net54),
    .A2(clknet_1_0__leaf_net899),
    .B1_N(net922),
    .X(net171));
 sky130_fd_sc_hd__a21bo_1 c249 (.A1(net170),
    .A2(net868),
    .B1_N(net702),
    .X(net172));
 sky130_fd_sc_hd__a31o_1 c250 (.A1(net25),
    .A2(net168),
    .A3(net788),
    .B1(net897),
    .X(net885));
 sky130_fd_sc_hd__sdfbbn_1 c251 (.CLK_N(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net171),
    .RESET_B(net169),
    .SCD(net871),
    .SCE(clknet_1_0__leaf_net899),
    .SET_B(net702),
    .Q(net174),
    .Q_N(net173));
 sky130_fd_sc_hd__a31o_1 c252 (.A1(net172),
    .A2(net169),
    .A3(net839),
    .B1(net151),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c253 (.A1(net175),
    .A2(net25),
    .B1_N(net64),
    .X(net176));
 sky130_fd_sc_hd__a21bo_1 c254 (.A1(net53),
    .A2(net173),
    .B1_N(net878),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 c255 (.A(net778),
    .X(net178));
 sky130_fd_sc_hd__a41o_1 c256 (.A1(net176),
    .A2(net55),
    .A3(net25),
    .A4(clknet_1_0__leaf_net899),
    .B1(net871),
    .X(net179));
 sky130_fd_sc_hd__a21bo_1 c257 (.A1(net174),
    .A2(net839),
    .B1_N(net907),
    .X(net852));
 sky130_fd_sc_hd__a21bo_1 c258 (.A1(net178),
    .A2(net169),
    .B1_N(net852),
    .X(net858));
 sky130_fd_sc_hd__a41o_1 c259 (.A1(net167),
    .A2(net174),
    .A3(clknet_1_0__leaf_net171),
    .A4(net868),
    .B1(net893),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net49),
    .A1(net149),
    .A2(net173),
    .A3(net150),
    .S0(net896),
    .S1(net852),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net181),
    .A1(clknet_1_0__leaf_net899),
    .A2(net173),
    .A3(net168),
    .S0(net656),
    .S1(net673),
    .X(net182));
 sky130_fd_sc_hd__a41o_1 c262 (.A1(clknet_1_1__leaf_net182),
    .A2(net174),
    .A3(net54),
    .A4(net169),
    .B1(net868),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net28),
    .A1(net181),
    .A2(clknet_1_0__leaf_net182),
    .A3(net54),
    .S0(net885),
    .S1(net168),
    .X(net184));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net842),
    .B(net73),
    .Y(net185));
 sky130_fd_sc_hd__xnor2_2 c265 (.A(net632),
    .B(net78),
    .Y(net186));
 sky130_fd_sc_hd__xnor2_1 c266 (.A(net185),
    .B(net73),
    .Y(net187));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net787),
    .A2(net186),
    .B1_N(net925),
    .X(net188));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net62),
    .B(net925),
    .Y(net189));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net185),
    .B(net927),
    .Y(net190));
 sky130_fd_sc_hd__a21bo_1 c270 (.A1(net846),
    .A2(net190),
    .B1_N(net927),
    .X(net191));
 sky130_fd_sc_hd__a21bo_2 c271 (.A1(net188),
    .A2(net190),
    .B1_N(net925),
    .X(net192));
 sky130_fd_sc_hd__a41o_1 c272 (.A1(net921),
    .A2(net65),
    .A3(net192),
    .A4(net925),
    .B1(net61),
    .X(net193));
 sky130_fd_sc_hd__a31o_2 c273 (.A1(net192),
    .A2(net189),
    .A3(net921),
    .B1(net925),
    .X(net194));
 sky130_fd_sc_hd__a31o_2 c274 (.A1(net190),
    .A2(net186),
    .A3(net789),
    .B1(net925),
    .X(net886));
 sky130_fd_sc_hd__a31o_2 c275 (.A1(net925),
    .A2(net787),
    .A3(net61),
    .B1(net192),
    .X(net195));
 sky130_fd_sc_hd__a21bo_1 c276 (.A1(net185),
    .A2(net886),
    .B1_N(net927),
    .X(net196));
 sky130_fd_sc_hd__a21bo_1 c277 (.A1(net195),
    .A2(net189),
    .B1_N(net193),
    .X(net197));
 sky130_fd_sc_hd__a21bo_1 c278 (.A1(net194),
    .A2(net886),
    .B1_N(net927),
    .X(net198));
 sky130_fd_sc_hd__mux4_2 c279 (.A0(net197),
    .A1(net198),
    .A2(net886),
    .A3(net188),
    .S0(net925),
    .S1(net921),
    .X(net199));
 sky130_fd_sc_hd__a41o_2 c280 (.A1(net886),
    .A2(net193),
    .A3(net921),
    .A4(net199),
    .B1(net925),
    .X(net200));
 sky130_fd_sc_hd__mux4_2 c281 (.A0(net200),
    .A1(net192),
    .A2(net199),
    .A3(net197),
    .S0(net189),
    .S1(net886),
    .X(net201));
 sky130_fd_sc_hd__a31o_4 c282 (.A1(net201),
    .A2(net192),
    .A3(net199),
    .B1(net925),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net196),
    .A1(net186),
    .A2(net201),
    .A3(net886),
    .S0(net189),
    .S1(net200),
    .X(net203));
 sky130_fd_sc_hd__mux4_2 c284 (.A0(net199),
    .A1(net203),
    .A2(net200),
    .A3(net188),
    .S0(net886),
    .S1(net921),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net203),
    .A1(net80),
    .A2(net204),
    .A3(net800),
    .S0(net192),
    .S1(net201),
    .X(net205));
 sky130_fd_sc_hd__a21bo_1 c286 (.A1(net98),
    .A2(net94),
    .B1_N(net926),
    .X(net206));
 sky130_fd_sc_hd__a21bo_1 c287 (.A1(net797),
    .A2(net98),
    .B1_N(net199),
    .X(net207));
 sky130_fd_sc_hd__a21bo_1 c288 (.A1(net68),
    .A2(net194),
    .B1_N(net78),
    .X(net208));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net831),
    .A2(net66),
    .B1_N(net916),
    .X(net209));
 sky130_fd_sc_hd__a31o_2 c290 (.A1(net208),
    .A2(net202),
    .A3(net98),
    .B1(net926),
    .X(net210));
 sky130_fd_sc_hd__a21bo_2 c291 (.A1(net209),
    .A2(net202),
    .B1_N(net206),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net821),
    .A1(net74),
    .A2(net192),
    .A3(net210),
    .S0(net186),
    .S1(net926),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net100),
    .A1(net68),
    .A2(net186),
    .A3(net211),
    .S0(net210),
    .S1(net976),
    .X(net213));
 sky130_fd_sc_hd__a21bo_1 c294 (.A1(net197),
    .A2(net97),
    .B1_N(net703),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net206),
    .A1(net210),
    .A2(net804),
    .A3(net68),
    .S0(net926),
    .S1(net916),
    .X(net215));
 sky130_fd_sc_hd__a21bo_1 c296 (.A1(net94),
    .A2(net100),
    .B1_N(net698),
    .X(net216));
 sky130_fd_sc_hd__buf_1 c297 (.A(net699),
    .X(net217));
 sky130_fd_sc_hd__a21bo_4 c298 (.A1(net61),
    .A2(net206),
    .B1_N(net804),
    .X(net218));
 sky130_fd_sc_hd__a21bo_4 c299 (.A1(net193),
    .A2(net209),
    .B1_N(net194),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 c300 (.A(net699),
    .X(net220));
 sky130_fd_sc_hd__a21bo_2 c301 (.A1(net220),
    .A2(net219),
    .B1_N(net698),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net186),
    .A1(net214),
    .A2(net821),
    .A3(net817),
    .S0(net80),
    .S1(net219),
    .X(net222));
 sky130_fd_sc_hd__sdfrtn_1 c303 (.CLK_N(clknet_4_5_0_clk),
    .D(net220),
    .RESET_B(net206),
    .SCD(net221),
    .SCE(net218),
    .Q(net223));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net216),
    .A1(net220),
    .A2(net221),
    .A3(net193),
    .S0(net219),
    .S1(net703),
    .X(net224));
 sky130_fd_sc_hd__a21bo_1 c305 (.A1(net188),
    .A2(net222),
    .B1_N(net805),
    .X(net225));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net225),
    .A2(net221),
    .A3(net223),
    .A4(net211),
    .B1(net926),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net222),
    .A1(net218),
    .A2(net225),
    .A3(net98),
    .S0(net223),
    .S1(net961),
    .X(net227));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net200),
    .B(net811),
    .Y(net228));
 sky130_fd_sc_hd__a21bo_2 c309 (.A1(net121),
    .A2(net83),
    .B1_N(net112),
    .X(net229));
 sky130_fd_sc_hd__a21bo_1 c310 (.A1(net93),
    .A2(net121),
    .B1_N(net817),
    .X(net230));
 sky130_fd_sc_hd__xnor2_1 c311 (.A(net817),
    .B(net698),
    .Y(net231));
 sky130_fd_sc_hd__xnor2_1 c312 (.A(net230),
    .B(net231),
    .Y(net232));
 sky130_fd_sc_hd__buf_1 c313 (.A(net695),
    .X(net233));
 sky130_fd_sc_hd__xnor2_4 c314 (.A(net836),
    .B(net93),
    .Y(net848));
 sky130_fd_sc_hd__a21bo_2 c315 (.A1(net843),
    .A2(net229),
    .B1_N(net909),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 c316 (.A(net970),
    .X(net235));
 sky130_fd_sc_hd__sdfrtp_4 c317 (.CLK(clknet_4_5_0_clk),
    .D(net202),
    .RESET_B(net204),
    .SCD(net229),
    .SCE(net699),
    .Q(net236));
 sky130_fd_sc_hd__a21bo_1 c318 (.A1(net78),
    .A2(net119),
    .B1_N(net928),
    .X(net237));
 sky130_fd_sc_hd__mux4_2 c319 (.A0(net121),
    .A1(net86),
    .A2(net73),
    .A3(net832),
    .S0(net926),
    .S1(net703),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 c320 (.A(net680),
    .X(net239));
 sky130_fd_sc_hd__buf_1 c321 (.A(net680),
    .X(net240));
 sky130_fd_sc_hd__a41o_1 c322 (.A1(net237),
    .A2(net909),
    .A3(net121),
    .A4(net238),
    .B1(net233),
    .X(net241));
 sky130_fd_sc_hd__a31o_1 c323 (.A1(net231),
    .A2(net233),
    .A3(net218),
    .B1(net240),
    .X(net242));
 sky130_fd_sc_hd__buf_1 c324 (.A(clknet_1_1__leaf_net782),
    .X(net243));
 sky130_fd_sc_hd__sdfbbn_2 c325 (.CLK_N(clknet_4_7_0_clk),
    .D(net210),
    .RESET_B(net969),
    .SCD(net235),
    .SCE(net240),
    .SET_B(net229),
    .Q(net876),
    .Q_N(net244));
 sky130_fd_sc_hd__sdfbbp_1 c326 (.CLK(clknet_4_5_0_clk),
    .D(net235),
    .RESET_B(net231),
    .SCD(clknet_1_0__leaf_net243),
    .SCE(net204),
    .SET_B(net228),
    .Q(net246),
    .Q_N(net245));
 sky130_fd_sc_hd__a21bo_2 c327 (.A1(net116),
    .A2(net240),
    .B1_N(net244),
    .X(net247));
 sky130_fd_sc_hd__a31o_1 c328 (.A1(net239),
    .A2(net237),
    .A3(net247),
    .B1(net238),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net86),
    .A1(net247),
    .A2(net200),
    .A3(net66),
    .S0(net229),
    .S1(net703),
    .X(net249));
 sky130_fd_sc_hd__sdfrtp_4 c330 (.CLK(clknet_4_7_0_clk),
    .D(net832),
    .RESET_B(net78),
    .SCD(net142),
    .SCE(net704),
    .Q(net250));
 sky130_fd_sc_hd__sdfrtp_2 c331 (.CLK(clknet_4_13_0_clk),
    .D(net119),
    .RESET_B(net958),
    .SCD(net922),
    .SCE(net142),
    .Q(net251));
 sky130_fd_sc_hd__clkbuf_1 c332 (.A(net776),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 c333 (.A(net775),
    .X(net872));
 sky130_fd_sc_hd__sdfsbp_1 c334 (.CLK(clknet_4_13_0_clk),
    .D(net130),
    .SCD(net973),
    .SCE(net142),
    .SET_B(net202),
    .Q(net882),
    .Q_N(net253));
 sky130_fd_sc_hd__clkbuf_1 c335 (.A(net695),
    .X(net254));
 sky130_fd_sc_hd__a31o_1 c336 (.A1(net249),
    .A2(net254),
    .A3(net872),
    .B1(net234),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c337 (.A1(net240),
    .A2(net909),
    .A3(net130),
    .A4(net250),
    .B1(net832),
    .X(net256));
 sky130_fd_sc_hd__a21bo_1 c338 (.A1(clknet_1_0__leaf_net243),
    .A2(net251),
    .B1_N(net119),
    .X(net257));
 sky130_fd_sc_hd__buf_1 c339 (.A(net784),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 c340 (.A(net786),
    .X(net259));
 sky130_fd_sc_hd__sdfsbp_1 c341 (.CLK(clknet_4_7_0_clk),
    .D(net254),
    .SCD(clknet_1_1__leaf_net243),
    .SCE(net256),
    .SET_B(net211),
    .Q(net877),
    .Q_N(net260));
 sky130_fd_sc_hd__a31o_2 c342 (.A1(net256),
    .A2(net843),
    .A3(net877),
    .B1(net872),
    .X(net261));
 sky130_fd_sc_hd__a31o_1 c343 (.A1(net107),
    .A2(clknet_1_1__leaf_net257),
    .A3(net261),
    .B1(net928),
    .X(net262));
 sky130_fd_sc_hd__a41o_1 c344 (.A1(clknet_1_0__leaf_net257),
    .A2(net90),
    .A3(net261),
    .A4(clknet_1_0__leaf_net262),
    .B1(net234),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net876),
    .A1(net130),
    .A2(net877),
    .A3(net138),
    .S0(clknet_1_0__leaf_net262),
    .S1(net698),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net19),
    .A1(clknet_1_1__leaf_net262),
    .A2(net877),
    .A3(net872),
    .S0(net674),
    .S1(net698),
    .X(net265));
 sky130_fd_sc_hd__sdfbbn_1 c347 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net265),
    .RESET_B(net219),
    .SCD(net261),
    .SCE(net882),
    .SET_B(net229),
    .Q(net267),
    .Q_N(net266));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(clknet_1_0__leaf_net262),
    .A1(net122),
    .A2(clknet_1_1__leaf_net265),
    .A3(net260),
    .S0(net251),
    .S1(net253),
    .X(net268));
 sky130_fd_sc_hd__a31o_1 c349 (.A1(net259),
    .A2(clknet_1_1__leaf_net262),
    .A3(net130),
    .B1(net675),
    .X(net892));
 sky130_fd_sc_hd__a41o_1 c350 (.A1(net23),
    .A2(net122),
    .A3(clknet_1_1__leaf_net262),
    .A4(net251),
    .B1(net266),
    .X(net269));
 sky130_fd_sc_hd__a41o_1 c351 (.A1(clknet_1_0__leaf_net269),
    .A2(net251),
    .A3(clknet_1_0__leaf_net892),
    .A4(net234),
    .B1(net252),
    .X(net270));
 sky130_fd_sc_hd__a21bo_1 c352 (.A1(net156),
    .A2(net154),
    .B1_N(net796),
    .X(net271));
 sky130_fd_sc_hd__buf_1 c353 (.A(net962),
    .X(net891));
 sky130_fd_sc_hd__xnor2_1 c354 (.A(net148),
    .B(net946),
    .Y(net272));
 sky130_fd_sc_hd__a31o_1 c355 (.A1(net73),
    .A2(net258),
    .A3(net271),
    .B1(net941),
    .X(net273));
 sky130_fd_sc_hd__a21bo_2 c356 (.A1(net153),
    .A2(net882),
    .B1_N(net32),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net128),
    .A1(net271),
    .A2(net32),
    .A3(net839),
    .S0(net274),
    .S1(net211),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net271),
    .A1(net148),
    .A2(net234),
    .A3(net274),
    .S0(clknet_1_0__leaf_net269),
    .S1(net662),
    .X(net276));
 sky130_fd_sc_hd__a21bo_1 c359 (.A1(net789),
    .A2(net155),
    .B1_N(net670),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 c360 (.A(net962),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 c361 (.A(net646),
    .X(net865));
 sky130_fd_sc_hd__buf_1 c362 (.A(net645),
    .X(net279));
 sky130_fd_sc_hd__a31o_1 c363 (.A1(net278),
    .A2(net163),
    .A3(net978),
    .B1(net904),
    .X(net884));
 sky130_fd_sc_hd__buf_1 c364 (.A(net779),
    .X(net280));
 sky130_fd_sc_hd__xnor2_1 c365 (.A(net154),
    .B(net73),
    .Y(net281));
 sky130_fd_sc_hd__buf_1 c366 (.A(clknet_1_1__leaf_net692),
    .X(net873));
 sky130_fd_sc_hd__a21bo_1 c367 (.A1(net155),
    .A2(net202),
    .B1_N(net670),
    .X(net282));
 sky130_fd_sc_hd__a21bo_1 c368 (.A1(net280),
    .A2(net157),
    .B1_N(net120),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 c369 (.A(net783),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 c370 (.A(net779),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 c371 (.A(net975),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net284),
    .A1(net278),
    .A2(net285),
    .A3(net274),
    .S0(net937),
    .S1(net891),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net285),
    .A1(clknet_1_1__leaf_net269),
    .A2(net155),
    .A3(net166),
    .S0(net281),
    .S1(net260),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net120),
    .A1(clknet_1_1__leaf_net269),
    .A2(net895),
    .A3(net128),
    .S0(net885),
    .S1(net863),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net277),
    .A1(net280),
    .A2(clknet_1_0__leaf_net873),
    .A3(net895),
    .S0(net888),
    .S1(clknet_1_0__leaf_net854),
    .X(net894));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net150),
    .A1(net181),
    .A2(net946),
    .A3(clknet_1_0__leaf_net894),
    .S0(net848),
    .S1(clknet_1_0__leaf_net854),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net149),
    .A1(net896),
    .A2(clknet_1_0__leaf_net894),
    .S0(net691),
    .S1(clknet_1_1__leaf_net854),
    .X(net290));
 sky130_fd_sc_hd__xnor2_2 c396 (.A(net79),
    .B(net74),
    .Y(net291));
 sky130_fd_sc_hd__xnor2_2 c397 (.A(net797),
    .B(net291),
    .Y(net292));
 sky130_fd_sc_hd__xnor2_4 c398 (.A(net931),
    .B(net699),
    .Y(net293));
 sky130_fd_sc_hd__xnor2_1 c399 (.A(net77),
    .B(net915),
    .Y(net294));
 sky130_fd_sc_hd__a31o_2 c400 (.A1(net919),
    .A2(net842),
    .A3(net293),
    .B1(net927),
    .X(net295));
 sky130_fd_sc_hd__xnor2_4 c401 (.A(net189),
    .B(net699),
    .Y(net296));
 sky130_fd_sc_hd__xnor2_4 c402 (.A(net915),
    .B(net919),
    .Y(net297));
 sky130_fd_sc_hd__a21bo_1 c403 (.A1(net845),
    .A2(net74),
    .B1_N(net296),
    .X(net869));
 sky130_fd_sc_hd__a21bo_2 c404 (.A1(net65),
    .A2(net295),
    .B1_N(net921),
    .X(net298));
 sky130_fd_sc_hd__xnor2_2 c405 (.A(net297),
    .B(net296),
    .Y(net299));
 sky130_fd_sc_hd__a41o_4 c406 (.A1(net299),
    .A2(net298),
    .A3(net293),
    .A4(net185),
    .B1(net927),
    .X(net300));
 sky130_fd_sc_hd__xnor2_2 c407 (.A(net298),
    .B(net920),
    .Y(net301));
 sky130_fd_sc_hd__a21bo_1 c408 (.A1(net294),
    .A2(net196),
    .B1_N(net924),
    .X(net302));
 sky130_fd_sc_hd__xnor2_4 c409 (.A(net190),
    .B(net297),
    .Y(net303));
 sky130_fd_sc_hd__xnor2_4 c410 (.A(net919),
    .B(net303),
    .Y(net304));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(net293),
    .A2(net301),
    .B1_N(net298),
    .X(net305));
 sky130_fd_sc_hd__xnor2_1 c412 (.A(net300),
    .B(net304),
    .Y(net306));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net304),
    .A2(net300),
    .B1_N(net306),
    .X(net307));
 sky130_fd_sc_hd__a21bo_1 c414 (.A1(net307),
    .A2(net304),
    .B1_N(net306),
    .X(net308));
 sky130_fd_sc_hd__xnor2_2 c415 (.A(net798),
    .B(net800),
    .Y(net309));
 sky130_fd_sc_hd__mux4_2 c416 (.A0(net305),
    .A1(net309),
    .A2(net308),
    .A3(net298),
    .S0(net915),
    .S1(net927),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net310),
    .A1(net198),
    .A2(net295),
    .A3(net308),
    .S0(net77),
    .S1(net305),
    .X(net311));
 sky130_fd_sc_hd__a21bo_2 c418 (.A1(net74),
    .A2(net194),
    .B1_N(net903),
    .X(net312));
 sky130_fd_sc_hd__a21bo_1 c419 (.A1(net306),
    .A2(net307),
    .B1_N(net219),
    .X(net313));
 sky130_fd_sc_hd__a21bo_4 c420 (.A1(net308),
    .A2(net846),
    .B1_N(net217),
    .X(net901));
 sky130_fd_sc_hd__a21bo_1 c421 (.A1(net214),
    .A2(net221),
    .B1_N(net313),
    .X(net314));
 sky130_fd_sc_hd__a21bo_2 c422 (.A1(net192),
    .A2(net917),
    .B1_N(net185),
    .X(net315));
 sky130_fd_sc_hd__a21bo_1 c423 (.A1(net314),
    .A2(net97),
    .B1_N(net214),
    .X(net316));
 sky130_fd_sc_hd__xnor2_2 c424 (.A(net315),
    .B(net303),
    .Y(net317));
 sky130_fd_sc_hd__xnor2_1 c425 (.A(net97),
    .B(net310),
    .Y(net318));
 sky130_fd_sc_hd__xnor2_1 c426 (.A(net318),
    .B(net298),
    .Y(net319));
 sky130_fd_sc_hd__a21bo_1 c427 (.A1(net313),
    .A2(net317),
    .B1_N(net307),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net301),
    .A1(net315),
    .A2(net318),
    .A3(net194),
    .S0(net312),
    .S1(net929),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 c429 (.A(net668),
    .X(net322));
 sky130_fd_sc_hd__a21bo_1 c430 (.A1(net207),
    .A2(net301),
    .B1_N(net668),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net298),
    .A1(net191),
    .A2(net317),
    .A3(net323),
    .S0(net312),
    .S1(net316),
    .X(net324));
 sky130_fd_sc_hd__a21bo_4 c432 (.A1(net845),
    .A2(net83),
    .B1_N(net668),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net194),
    .A1(net920),
    .A2(net314),
    .A3(net301),
    .S0(net317),
    .S1(net312),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 c434 (.A(net668),
    .X(net327));
 sky130_fd_sc_hd__a21bo_1 c435 (.A1(net207),
    .A2(net308),
    .B1_N(clknet_1_1__leaf_net706),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net317),
    .A1(net323),
    .A2(net327),
    .A3(net77),
    .S0(net320),
    .S1(clknet_1_1__leaf_net706),
    .X(net329));
 sky130_fd_sc_hd__a21bo_1 c437 (.A1(net804),
    .A2(net223),
    .B1_N(net325),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net328),
    .A1(net305),
    .A2(net808),
    .A3(net191),
    .S0(net301),
    .S1(net709),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net320),
    .A1(net314),
    .A2(net313),
    .A3(net307),
    .S0(net310),
    .S1(net711),
    .X(net332));
 sky130_fd_sc_hd__sdfstp_1 c440 (.CLK(clknet_4_7_0_clk),
    .D(net248),
    .SCD(net316),
    .SCE(net123),
    .SET_B(net961),
    .Q(net333));
 sky130_fd_sc_hd__xnor2_2 c441 (.A(net325),
    .B(net699),
    .Y(net334));
 sky130_fd_sc_hd__buf_1 c442 (.A(net690),
    .X(net335));
 sky130_fd_sc_hd__xnor2_1 c443 (.A(net247),
    .B(net295),
    .Y(net336));
 sky130_fd_sc_hd__xnor2_2 c444 (.A(net334),
    .B(net79),
    .Y(net337));
 sky130_fd_sc_hd__a31o_2 c445 (.A1(net303),
    .A2(net337),
    .A3(net335),
    .B1(net245),
    .X(net338));
 sky130_fd_sc_hd__xnor2_1 c446 (.A(net338),
    .B(net711),
    .Y(net339));
 sky130_fd_sc_hd__xnor2_1 c447 (.A(net337),
    .B(net338),
    .Y(net340));
 sky130_fd_sc_hd__dlymetal6s2s_1 c448 (.A(net690),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net340),
    .A1(net791),
    .A2(net334),
    .A3(net303),
    .S0(net704),
    .S1(net710),
    .X(net342));
 sky130_fd_sc_hd__xnor2_1 c450 (.A(net837),
    .B(net336),
    .Y(net343));
 sky130_fd_sc_hd__a41o_1 c451 (.A1(net217),
    .A2(net337),
    .A3(net341),
    .A4(net330),
    .B1(net340),
    .X(net344));
 sky130_fd_sc_hd__xnor2_1 c452 (.A(net295),
    .B(net246),
    .Y(net345));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(net339),
    .A1(net312),
    .A2(net837),
    .A3(net247),
    .S0(net911),
    .S1(net337),
    .X(net346));
 sky130_fd_sc_hd__a21bo_1 c454 (.A1(net342),
    .A2(net339),
    .B1_N(net911),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net336),
    .A1(net293),
    .A2(net322),
    .A3(net312),
    .S0(net911),
    .S1(net303),
    .X(net348));
 sky130_fd_sc_hd__sdfstp_2 c456 (.CLK(clknet_4_6_0_clk),
    .D(net817),
    .SCD(net335),
    .SCE(net911),
    .SET_B(net123),
    .Q(net859));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net241),
    .A1(net110),
    .A2(net337),
    .A3(net333),
    .S0(net247),
    .S1(net714),
    .X(net349));
 sky130_fd_sc_hd__a41o_1 c458 (.A1(net246),
    .A2(net903),
    .A3(net911),
    .A4(net714),
    .B1(net715),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net350),
    .A1(net347),
    .A2(net295),
    .A3(net303),
    .S0(net911),
    .S1(net714),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net247),
    .A1(net350),
    .A2(net859),
    .A3(net911),
    .S1(net715),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net342),
    .A1(net350),
    .A2(net315),
    .A3(net303),
    .S0(net667),
    .S1(net714),
    .X(net353));
 sky130_fd_sc_hd__a31o_1 c462 (.A1(net344),
    .A2(net202),
    .A3(net920),
    .B1(net911),
    .X(net354));
 sky130_fd_sc_hd__a31o_1 c463 (.A1(net138),
    .A2(net876),
    .A3(net928),
    .B1(net913),
    .X(net355));
 sky130_fd_sc_hd__buf_1 c464 (.A(net774),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 c465 (.A(net773),
    .X(net357));
 sky130_fd_sc_hd__buf_1 c466 (.A(clknet_1_0__leaf_net692),
    .X(net861));
 sky130_fd_sc_hd__a31o_1 c467 (.A1(net811),
    .A2(net106),
    .A3(net912),
    .B1(net705),
    .X(net358));
 sky130_fd_sc_hd__a21bo_1 c468 (.A1(net937),
    .A2(net920),
    .B1_N(net843),
    .X(net359));
 sky130_fd_sc_hd__a21bo_1 c469 (.A1(net856),
    .A2(net356),
    .B1_N(net659),
    .X(net360));
 sky130_fd_sc_hd__buf_1 c470 (.A(clknet_1_1__leaf_net692),
    .X(net860));
 sky130_fd_sc_hd__buf_1 c471 (.A(clknet_1_0__leaf_net692),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(clknet_1_0__leaf_net361),
    .A1(net335),
    .A2(clknet_1_0__leaf_net861),
    .A3(net250),
    .S0(net705),
    .S1(net715),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net928),
    .A1(clknet_1_1__leaf_net362),
    .A2(net360),
    .A3(net920),
    .S0(net260),
    .S1(net696),
    .X(net363));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(net335),
    .A2(net344),
    .B1_N(clknet_1_0__leaf_net861),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 c475 (.A(net687),
    .X(net857));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net843),
    .A1(clknet_1_0__leaf_net860),
    .A2(net932),
    .A3(net913),
    .S0(net928),
    .S1(net716),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net219),
    .A1(clknet_1_1__leaf_net361),
    .A2(clknet_1_1__leaf_net364),
    .A3(net920),
    .S0(net928),
    .S1(net716),
    .X(net366));
 sky130_fd_sc_hd__a31o_1 c478 (.A1(net366),
    .A2(net920),
    .A3(net932),
    .B1(net716),
    .X(net367));
 sky130_fd_sc_hd__a31o_1 c479 (.A1(net330),
    .A2(clknet_1_0__leaf_net860),
    .A3(clknet_1_1__leaf_net362),
    .B1(net932),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net368),
    .A1(net360),
    .A2(net138),
    .A3(net843),
    .S0(net259),
    .S1(clknet_1_1__leaf_net364),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net360),
    .A1(clknet_1_1__leaf_net362),
    .A2(net259),
    .A3(net358),
    .S0(net716),
    .S1(net717),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net358),
    .A1(clknet_1_1__leaf_net362),
    .A2(net219),
    .A3(net359),
    .S0(net715),
    .S1(net716),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net920),
    .A1(net219),
    .A2(clknet_1_0__leaf_net371),
    .A3(clknet_1_1__leaf_net367),
    .S0(clknet_1_0__leaf_net861),
    .S1(net717),
    .X(net372));
 sky130_fd_sc_hd__a41o_1 c484 (.A1(net922),
    .A2(net978),
    .A3(net272),
    .A4(net274),
    .B1(net957),
    .X(net373));
 sky130_fd_sc_hd__a31o_2 c485 (.A1(net77),
    .A2(net135),
    .A3(net859),
    .B1(net937),
    .X(net374));
 sky130_fd_sc_hd__a41o_1 c486 (.A1(net850),
    .A2(clknet_1_0__leaf_net873),
    .A3(net112),
    .A4(net662),
    .B1(net666),
    .X(net375));
 sky130_fd_sc_hd__a31o_1 c487 (.A1(net112),
    .A2(net922),
    .A3(net920),
    .B1(net850),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net365),
    .A1(net376),
    .A2(net904),
    .A3(net909),
    .S0(net356),
    .S1(net689),
    .X(net377));
 sky130_fd_sc_hd__a41o_1 c489 (.A1(net356),
    .A2(net202),
    .A3(clknet_1_0__leaf_net860),
    .A4(net244),
    .B1(net805),
    .X(net862));
 sky130_fd_sc_hd__sdfstp_1 c490 (.CLK(clknet_4_14_0_clk),
    .D(net166),
    .SCD(net953),
    .SCE(clknet_1_0__leaf_net862),
    .SET_B(clknet_1_0__leaf_net873),
    .Q(net378));
 sky130_fd_sc_hd__a41o_1 c491 (.A1(clknet_1_0__leaf_net377),
    .A2(net378),
    .A3(net112),
    .A4(net32),
    .B1(net376),
    .X(net379));
 sky130_fd_sc_hd__sdfbbn_1 c492 (.CLK_N(clknet_4_12_0_clk),
    .D(net791),
    .RESET_B(net974),
    .SCD(net922),
    .SCE(clknet_1_0__leaf_net862),
    .SET_B(net965),
    .Q(net380));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net856),
    .A1(net941),
    .A2(clknet_1_0__leaf_net862),
    .A3(net274),
    .S0(clknet_1_1__leaf_net377),
    .S1(net694),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net380),
    .A1(net932),
    .A2(net279),
    .A3(clknet_1_0__leaf_net862),
    .S0(net942),
    .S1(net953),
    .X(net382));
 sky130_fd_sc_hd__a41o_1 c495 (.A1(net792),
    .A2(net378),
    .A3(net374),
    .A4(net689),
    .B1(net718),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net374),
    .A1(net378),
    .A2(net811),
    .A3(clknet_1_0__leaf_net860),
    .S0(clknet_1_0__leaf_net861),
    .S1(net707),
    .X(net384));
 sky130_fd_sc_hd__sdfbbp_1 c497 (.CLK(clknet_4_14_0_clk),
    .D(net375),
    .RESET_B(clknet_1_0__leaf_net862),
    .SCD(net32),
    .SCE(clknet_1_0__leaf_net860),
    .SET_B(net950),
    .Q(net385));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net202),
    .A1(net918),
    .A2(clknet_1_1__leaf_net862),
    .A3(net694),
    .S0(clknet_1_0__leaf_net874),
    .S1(net718),
    .X(net386));
 sky130_fd_sc_hd__sdfbbn_1 c499 (.CLK_N(clknet_4_12_0_clk),
    .D(net378),
    .RESET_B(net166),
    .SCD(net869),
    .SCE(net707),
    .SET_B(net719),
    .Q(net388),
    .Q_N(net387));
 sky130_fd_sc_hd__mux4_2 c500 (.A0(net388),
    .A1(net32),
    .A2(net941),
    .A3(net914),
    .S0(net662),
    .S1(net721),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net385),
    .A1(net389),
    .A2(net274),
    .A3(net978),
    .S0(net951),
    .S1(net721),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net804),
    .A1(net166),
    .A2(net378),
    .A3(net719),
    .S0(net721),
    .S1(net722),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net238),
    .A1(net376),
    .A2(net948),
    .A3(net387),
    .S0(net658),
    .S1(net721),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net274),
    .A1(net956),
    .A2(net374),
    .A3(net392),
    .S0(net691),
    .S1(net722),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net159),
    .A1(net376),
    .A2(net933),
    .A3(net866),
    .S0(net722),
    .S1(net723),
    .X(net394));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net931),
    .B(net929),
    .Y(net395));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net794),
    .B(net195),
    .Y(net396));
 sky130_fd_sc_hd__xnor2_2 c530 (.A(net800),
    .B(net299),
    .Y(net397));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net304),
    .B(net395),
    .Y(net398));
 sky130_fd_sc_hd__xnor2_1 c532 (.A(net398),
    .B(net397),
    .Y(net399));
 sky130_fd_sc_hd__a21bo_1 c533 (.A1(net399),
    .A2(net792),
    .B1_N(net398),
    .X(net400));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net296),
    .B(net931),
    .Y(net401));
 sky130_fd_sc_hd__mux4_2 c535 (.A0(net794),
    .A1(net296),
    .A2(net300),
    .A3(net401),
    .S0(net398),
    .S1(net395),
    .X(net402));
 sky130_fd_sc_hd__xnor2_1 c536 (.A(net299),
    .B(net311),
    .Y(net403));
 sky130_fd_sc_hd__a21bo_1 c537 (.A1(net402),
    .A2(net398),
    .B1_N(net924),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net400),
    .A1(net403),
    .A2(net302),
    .A3(net395),
    .S0(net398),
    .S1(net396),
    .X(net405));
 sky130_fd_sc_hd__a21bo_1 c539 (.A1(net294),
    .A2(net399),
    .B1_N(clknet_1_1__leaf_net724),
    .X(net406));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(clknet_1_1__leaf_net406),
    .A2(net398),
    .B1_N(net302),
    .X(net407));
 sky130_fd_sc_hd__a21bo_1 c541 (.A1(net302),
    .A2(net296),
    .B1_N(clknet_1_1__leaf_net724),
    .X(net408));
 sky130_fd_sc_hd__a41o_1 c542 (.A1(net397),
    .A2(net404),
    .A3(net399),
    .A4(net931),
    .B1(net699),
    .X(net409));
 sky130_fd_sc_hd__a21bo_1 c543 (.A1(net401),
    .A2(clknet_1_0__leaf_net407),
    .B1_N(net398),
    .X(net410));
 sky130_fd_sc_hd__a21bo_1 c544 (.A1(clknet_1_0__leaf_net410),
    .A2(net402),
    .B1_N(clknet_1_0__leaf_net407),
    .X(net411));
 sky130_fd_sc_hd__a41o_1 c545 (.A1(net395),
    .A2(net401),
    .A3(clknet_1_1__leaf_net410),
    .A4(clknet_1_0__leaf_net407),
    .B1(net402),
    .X(net412));
 sky130_fd_sc_hd__buf_2 c546 (.A(net663),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_1__leaf_net411),
    .A1(net413),
    .A2(clknet_1_0__leaf_net412),
    .A3(net404),
    .S0(clknet_1_0__leaf_net406),
    .S1(net296),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 c548 (.A(net663),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net409),
    .A1(net415),
    .A2(clknet_1_0__leaf_net410),
    .A3(net395),
    .S0(net402),
    .S1(net294),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_4 c550 (.A(net682),
    .X(net417));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net791),
    .A2(net901),
    .B1_N(net632),
    .X(net418));
 sky130_fd_sc_hd__a21bo_1 c552 (.A1(net297),
    .A2(clknet_1_0__leaf_net706),
    .B1_N(net709),
    .X(net419));
 sky130_fd_sc_hd__a31o_1 c553 (.A1(net309),
    .A2(net327),
    .A3(net901),
    .B1(net417),
    .X(net420));
 sky130_fd_sc_hd__buf_1 c554 (.A(clknet_1_1__leaf_net781),
    .X(net421));
 sky130_fd_sc_hd__a21bo_1 c555 (.A1(clknet_1_0__leaf_net421),
    .A2(net417),
    .B1_N(net710),
    .X(net422));
 sky130_fd_sc_hd__a21bo_1 c556 (.A1(net420),
    .A2(net921),
    .B1_N(clknet_1_1__leaf_net421),
    .X(net423));
 sky130_fd_sc_hd__mux4_2 c557 (.A0(net418),
    .A1(net901),
    .A2(net417),
    .A3(net921),
    .S0(net924),
    .S1(net710),
    .X(net424));
 sky130_fd_sc_hd__buf_1 c558 (.A(clknet_1_1__leaf_net780),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net682),
    .X(net426));
 sky130_fd_sc_hd__buf_1 c560 (.A(net682),
    .X(net427));
 sky130_fd_sc_hd__a21bo_1 c561 (.A1(net418),
    .A2(clknet_1_1__leaf_net425),
    .B1_N(clknet_1_0__leaf_net422),
    .X(net428));
 sky130_fd_sc_hd__sdfbbn_2 c562 (.CLK_N(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net425),
    .RESET_B(net325),
    .SCD(net83),
    .SCE(clknet_1_1__leaf_net421),
    .SET_B(clknet_1_0__leaf_net423),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__buf_2 c563 (.A(net682),
    .X(net889));
 sky130_fd_sc_hd__buf_1 c564 (.A(clknet_1_0__leaf_net780),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net420),
    .A1(net323),
    .A2(clknet_1_0__leaf_net431),
    .A3(clknet_1_1__leaf_net419),
    .S0(net327),
    .S1(net221),
    .X(net432));
 sky130_fd_sc_hd__buf_1 c566 (.A(clknet_1_0__leaf_net693),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_0__leaf_net433),
    .A1(net413),
    .A2(net403),
    .A3(net97),
    .S0(net223),
    .S1(clknet_1_1__leaf_net408),
    .X(net434));
 sky130_fd_sc_hd__a21bo_1 c568 (.A1(net846),
    .A2(clknet_1_0__leaf_net422),
    .B1_N(net726),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net632),
    .A1(net889),
    .A2(clknet_1_0__leaf_net425),
    .A3(net429),
    .S0(net725),
    .S1(net727),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(clknet_1_0__leaf_net431),
    .A1(clknet_1_0__leaf_net435),
    .A2(net915),
    .A3(clknet_1_1__leaf_net433),
    .S0(clknet_1_1__leaf_net425),
    .S1(net420),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(clknet_1_0__leaf_net435),
    .A1(net427),
    .A2(net426),
    .A3(net420),
    .S0(clknet_1_0__leaf_net437),
    .S1(net726),
    .X(net438));
 sky130_fd_sc_hd__a21bo_1 c572 (.A1(net83),
    .A2(net396),
    .B1_N(net927),
    .X(net439));
 sky130_fd_sc_hd__xnor2_1 c573 (.A(net338),
    .B(net713),
    .Y(net440));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net123),
    .A1(net903),
    .A2(clknet_1_1__leaf_net435),
    .A3(net343),
    .S0(clknet_1_1__leaf_net423),
    .S1(net417),
    .X(net441));
 sky130_fd_sc_hd__buf_1 c575 (.A(net697),
    .X(net442));
 sky130_fd_sc_hd__xnor2_1 c576 (.A(net315),
    .B(net831),
    .Y(net443));
 sky130_fd_sc_hd__clkbuf_1 c577 (.A(net785),
    .X(net444));
 sky130_fd_sc_hd__xnor2_2 c578 (.A(net440),
    .B(net338),
    .Y(net445));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net697),
    .X(net446));
 sky130_fd_sc_hd__xnor2_1 c580 (.A(clknet_1_1__leaf_net431),
    .B(net417),
    .Y(net447));
 sky130_fd_sc_hd__a21bo_1 c581 (.A1(net447),
    .A2(net859),
    .B1_N(net236),
    .X(net448));
 sky130_fd_sc_hd__buf_1 c582 (.A(clknet_1_0__leaf_net782),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 c583 (.A(net777),
    .X(net450));
 sky130_fd_sc_hd__a31o_1 c584 (.A1(net347),
    .A2(clknet_1_0__leaf_net407),
    .A3(clknet_1_1__leaf_net422),
    .B1(net923),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net448),
    .A1(net322),
    .A2(clknet_1_0__leaf_net416),
    .A3(clknet_1_1__leaf_net422),
    .S0(net911),
    .S1(net923),
    .X(net452));
 sky130_fd_sc_hd__xnor2_1 c586 (.A(net236),
    .B(net106),
    .Y(net453));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net450),
    .A1(clknet_1_0__leaf_net437),
    .A2(clknet_1_0__leaf_net422),
    .A3(net911),
    .S0(net709),
    .S1(net713),
    .X(net454));
 sky130_fd_sc_hd__a21bo_1 c588 (.A1(net236),
    .A2(clknet_1_1__leaf_net693),
    .B1_N(net935),
    .X(net849));
 sky130_fd_sc_hd__xnor2_1 c589 (.A(net445),
    .B(net417),
    .Y(net455));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net453),
    .A1(net455),
    .A2(clknet_1_0__leaf_net423),
    .A3(clknet_1_1__leaf_net449),
    .S0(net417),
    .S1(clknet_1_0__leaf_net416),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net444),
    .A1(net451),
    .A2(net325),
    .A3(net903),
    .S0(clknet_1_0__leaf_net407),
    .S1(net710),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net442),
    .A1(clknet_1_0__leaf_net457),
    .A2(net445),
    .A3(net713),
    .S0(net935),
    .S1(net851),
    .X(net458));
 sky130_fd_sc_hd__buf_1 c593 (.A(clknet_1_0__leaf_net781),
    .X(net459));
 sky130_fd_sc_hd__sdfbbp_1 c594 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net437),
    .RESET_B(net250),
    .SCD(net261),
    .SCE(net909),
    .SET_B(clknet_1_0__leaf_net364),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__a41o_1 c595 (.A1(net259),
    .A2(clknet_1_0__leaf_net364),
    .A3(net77),
    .A4(net937),
    .B1(net732),
    .X(net462));
 sky130_fd_sc_hd__sdfbbn_1 c596 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net428),
    .RESET_B(net972),
    .SCD(net912),
    .SCE(net923),
    .SET_B(net963),
    .Q(net464),
    .Q_N(net463));
 sky130_fd_sc_hd__sdfbbn_1 c597 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net372),
    .RESET_B(net461),
    .SCD(net856),
    .SCE(clknet_1_1__leaf_net407),
    .SET_B(net905),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__sedfxbp_2 c598 (.CLK(clknet_4_3_0_clk),
    .D(net343),
    .DE(net912),
    .SCD(clknet_1_1__leaf_net422),
    .SCE(net429),
    .Q(net468),
    .Q_N(net467));
 sky130_fd_sc_hd__sdfbbp_1 c599 (.CLK(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net428),
    .RESET_B(net971),
    .SCD(net396),
    .SCE(net359),
    .SET_B(net961),
    .Q(net470),
    .Q_N(net469));
 sky130_fd_sc_hd__mux4_2 c600 (.A0(net464),
    .A1(net465),
    .A2(net261),
    .A3(net469),
    .S0(net924),
    .S1(net791),
    .X(net471));
 sky130_fd_sc_hd__sdfbbn_2 c601 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net367),
    .RESET_B(clknet_1_0__leaf_net371),
    .SCD(clknet_1_1__leaf_net437),
    .SCE(net905),
    .SET_B(clknet_1_1__leaf_net407),
    .Q(net473),
    .Q_N(net472));
 sky130_fd_sc_hd__a41o_1 c602 (.A1(clknet_1_1__leaf_net422),
    .A2(clknet_1_0__leaf_net407),
    .A3(net463),
    .A4(net708),
    .B1(net732),
    .X(net474));
 sky130_fd_sc_hd__a41o_1 c603 (.A1(net359),
    .A2(net462),
    .A3(net470),
    .A4(net267),
    .B1(net905),
    .X(net475));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_4_6_0_clk),
    .D(net417),
    .RESET_B(net967),
    .SCD(net471),
    .SCE(clknet_1_0__leaf_net372),
    .SET_B(net932),
    .Q(net477),
    .Q_N(net476));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_0__leaf_net364),
    .A1(net889),
    .A2(net463),
    .A3(net918),
    .S0(clknet_1_1__leaf_net428),
    .S1(net261),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net808),
    .A1(clknet_1_0__leaf_net474),
    .A2(net912),
    .A3(net476),
    .S0(net704),
    .S1(net880),
    .X(net479));
 sky130_fd_sc_hd__a41o_1 c607 (.A1(clknet_1_0__leaf_net362),
    .A2(clknet_1_1__leaf_net860),
    .A3(net704),
    .A4(net712),
    .B1(net880),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net466),
    .A1(net915),
    .A2(clknet_1_0__leaf_net362),
    .A3(net463),
    .S0(net728),
    .S1(net880),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net480),
    .A1(clknet_1_1__leaf_net457),
    .A2(clknet_1_0__leaf_net474),
    .A3(clknet_1_0__leaf_net362),
    .S0(clknet_1_1__leaf_net479),
    .S1(net880),
    .X(net482));
 sky130_fd_sc_hd__a41o_1 c610 (.A1(net261),
    .A2(net464),
    .A3(clknet_1_1__leaf_net479),
    .A4(net905),
    .B1(net469),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net477),
    .A1(clknet_1_1__leaf_net479),
    .A2(net471),
    .A3(net472),
    .S0(net935),
    .S1(net880),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net466),
    .A1(net918),
    .A2(net461),
    .A3(net932),
    .S0(net880),
    .S1(net735),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net481),
    .A1(net485),
    .A2(clknet_1_1__leaf_net407),
    .A3(net359),
    .S0(net678),
    .S1(net734),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net485),
    .A1(clknet_1_0__leaf_net479),
    .A2(net460),
    .A3(net267),
    .S0(net733),
    .S1(net735),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net325),
    .A1(net475),
    .A2(net79),
    .A3(net913),
    .S0(net485),
    .S1(net471),
    .X(net488));
 sky130_fd_sc_hd__a41o_1 c616 (.A1(clknet_1_1__leaf_net407),
    .A2(net907),
    .A3(net856),
    .A4(net933),
    .B1(net721),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net446),
    .A1(net374),
    .A2(net471),
    .A3(net811),
    .S0(clknet_1_0__leaf_net860),
    .S1(net795),
    .X(net490));
 sky130_fd_sc_hd__a41o_1 c618 (.A1(clknet_1_1__leaf_net407),
    .A2(net473),
    .A3(net953),
    .A4(net266),
    .B1(net720),
    .X(net491));
 sky130_fd_sc_hd__sdfbbp_1 c619 (.CLK(clknet_4_9_0_clk),
    .D(net267),
    .RESET_B(clknet_1_0__leaf_net489),
    .SCD(clknet_1_1__leaf_net860),
    .SCE(clknet_1_0__leaf_net394),
    .SET_B(net471),
    .Q(net493),
    .Q_N(net492));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net827),
    .A1(net832),
    .A2(net838),
    .A3(net834),
    .S0(net830),
    .S1(net801),
    .X(net0));
 sky130_fd_sc_hd__sdfbbn_1 c620 (.CLK_N(clknet_4_11_0_clk),
    .D(net493),
    .RESET_B(net812),
    .SCD(net906),
    .SCE(clknet_1_0__leaf_net489),
    .SET_B(net966),
    .Q(net495),
    .Q_N(net494));
 sky130_fd_sc_hd__a41o_1 c621 (.A1(net471),
    .A2(net491),
    .A3(net909),
    .A4(net32),
    .B1(net949),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net495),
    .A1(net906),
    .A2(clknet_1_1__leaf_net860),
    .A3(net907),
    .S0(clknet_1_1__leaf_net693),
    .S1(net697),
    .X(net853));
 sky130_fd_sc_hd__a41o_1 c623 (.A1(net495),
    .A2(net799),
    .A3(clknet_1_1__leaf_net407),
    .A4(net953),
    .B1(net913),
    .X(net497));
 sky130_fd_sc_hd__a41o_1 c624 (.A1(clknet_1_1__leaf_net371),
    .A2(net497),
    .A3(net811),
    .A4(clknet_1_1__leaf_net860),
    .B1(net933),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net906),
    .A1(net374),
    .A2(net889),
    .A3(clknet_1_0__leaf_net394),
    .S0(net811),
    .S1(net494),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net272),
    .A1(clknet_1_1__leaf_net435),
    .A2(clknet_1_1__leaf_net489),
    .A3(net472),
    .S0(net953),
    .S1(net870),
    .X(net500));
 sky130_fd_sc_hd__a41o_1 c627 (.A1(net32),
    .A2(net496),
    .A3(net471),
    .A4(clknet_1_0__leaf_net860),
    .B1(net736),
    .X(net501));
 sky130_fd_sc_hd__a41o_1 c628 (.A1(net811),
    .A2(net468),
    .A3(net661),
    .A4(net721),
    .B1(net737),
    .X(net502));
 sky130_fd_sc_hd__sdfbbn_1 c629 (.CLK_N(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net407),
    .RESET_B(net498),
    .SCD(net32),
    .SCE(net870),
    .SET_B(net737),
    .Q(net503));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net814),
    .A1(net835),
    .A2(net834),
    .A3(net840),
    .S0(net836),
    .S1(net801),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net279),
    .A1(net937),
    .A2(net914),
    .A3(net661),
    .S0(net721),
    .S1(net736),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net443),
    .A1(clknet_1_0__leaf_net873),
    .A2(clknet_1_0__leaf_net377),
    .A3(net914),
    .S0(net870),
    .S1(net737),
    .X(net505));
 sky130_fd_sc_hd__a41o_1 c632 (.A1(net503),
    .A2(clknet_1_1__leaf_net861),
    .A3(net870),
    .A4(net737),
    .B1(net738),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net341),
    .A1(clknet_1_1__leaf_net394),
    .A2(net492),
    .A3(net721),
    .S0(net736),
    .S1(net738),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net506),
    .A1(clknet_1_1__leaf_net861),
    .A2(net374),
    .A3(net736),
    .S0(net738),
    .S1(net739),
    .X(net508));
 sky130_fd_sc_hd__a41o_1 c635 (.A1(net389),
    .A2(net736),
    .A3(net737),
    .A4(net738),
    .B1(net740),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net502),
    .A1(net504),
    .A2(net392),
    .A3(clknet_1_1__leaf_net394),
    .S0(net904),
    .S1(net738),
    .X(net510));
 sky130_fd_sc_hd__a41o_1 c637 (.A1(net509),
    .A2(net901),
    .A3(net728),
    .A4(net738),
    .B1(clknet_1_1__leaf_net741),
    .X(net511));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net828),
    .A1(net1),
    .A2(net826),
    .A3(net829),
    .S0(net3),
    .S1(net837),
    .X(net2));
 sky130_fd_sc_hd__a21bo_1 c65 (.A1(net801),
    .A2(net847),
    .B1_N(net814),
    .X(net3));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net0),
    .B(net825),
    .Y(net4));
 sky130_fd_sc_hd__xnor2_4 c660 (.A(net929),
    .B(net300),
    .Y(net512));
 sky130_fd_sc_hd__a31o_1 c661 (.A1(net300),
    .A2(net413),
    .A3(net663),
    .B1(clknet_1_0__leaf_net724),
    .X(net513));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net512),
    .B(net397),
    .Y(net514));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net195),
    .B(net514),
    .Y(net515));
 sky130_fd_sc_hd__xnor2_1 c664 (.A(net196),
    .B(clknet_1_1__leaf_net724),
    .Y(net516));
 sky130_fd_sc_hd__xnor2_1 c665 (.A(clknet_1_0__leaf_net513),
    .B(net794),
    .Y(net517));
 sky130_fd_sc_hd__a31o_1 c666 (.A1(net514),
    .A2(net903),
    .A3(clknet_1_1__leaf_net516),
    .B1(clknet_1_1__leaf_net513),
    .X(net518));
 sky130_fd_sc_hd__a21bo_1 c667 (.A1(clknet_1_1__leaf_net517),
    .A2(net924),
    .B1_N(net663),
    .X(net519));
 sky130_fd_sc_hd__xnor2_1 c668 (.A(clknet_1_0__leaf_net516),
    .B(clknet_1_1__leaf_net408),
    .Y(net520));
 sky130_fd_sc_hd__xnor2_1 c669 (.A(clknet_1_0__leaf_net520),
    .B(clknet_1_0__leaf_net724),
    .Y(net521));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net798),
    .B(net845),
    .Y(net5));
 sky130_fd_sc_hd__buf_1 c670 (.A(net664),
    .X(net522));
 sky130_fd_sc_hd__xnor2_4 c671 (.A(net512),
    .B(net699),
    .Y(net523));
 sky130_fd_sc_hd__xnor2_4 c672 (.A(net903),
    .B(net523),
    .Y(net524));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net198),
    .A1(net523),
    .A2(clknet_1_1__leaf_net518),
    .A3(net524),
    .S0(net514),
    .S1(net663),
    .X(net525));
 sky130_fd_sc_hd__xnor2_1 c674 (.A(net522),
    .B(clknet_1_0__leaf_net408),
    .Y(net526));
 sky130_fd_sc_hd__xnor2_2 c675 (.A(net398),
    .B(net915),
    .Y(net527));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(clknet_1_1__leaf_net520),
    .A1(net523),
    .A2(net522),
    .A3(net908),
    .S0(net663),
    .S1(net665),
    .X(net528));
 sky130_fd_sc_hd__xnor2_1 c677 (.A(clknet_1_0__leaf_net517),
    .B(net663),
    .Y(net529));
 sky130_fd_sc_hd__clkbuf_4 c678 (.A(net664),
    .X(net530));
 sky130_fd_sc_hd__xnor2_1 c679 (.A(clknet_1_0__leaf_net529),
    .B(net523),
    .Y(net531));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net4),
    .B(net807),
    .Y(net6));
 sky130_fd_sc_hd__buf_1 c680 (.A(clknet_1_0__leaf_net693),
    .X(net532));
 sky130_fd_sc_hd__sdfbbp_1 c681 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net528),
    .RESET_B(clknet_1_0__leaf_net531),
    .SCD(net524),
    .SCE(clknet_1_0__leaf_net529),
    .SET_B(net665),
    .Q(net534),
    .Q_N(net533));
 sky130_fd_sc_hd__a21bo_1 c682 (.A1(net185),
    .A2(clknet_1_1__leaf_net529),
    .B1_N(net429),
    .X(net535));
 sky130_fd_sc_hd__a31o_1 c683 (.A1(net427),
    .A2(net524),
    .A3(clknet_1_0__leaf_net535),
    .B1(net903),
    .X(net536));
 sky130_fd_sc_hd__a21bo_1 c684 (.A1(clknet_1_0__leaf_net532),
    .A2(clknet_1_1__leaf_net526),
    .B1_N(clknet_1_0__leaf_net529),
    .X(net537));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net921),
    .A2(clknet_1_0__leaf_net535),
    .A3(clknet_1_1__leaf_net537),
    .B1(net730),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(clknet_1_0__leaf_net436),
    .A1(clknet_1_0__leaf_net518),
    .A2(net929),
    .A3(clknet_1_0__leaf_net526),
    .S0(net97),
    .S1(clknet_1_0__leaf_net408),
    .X(net539));
 sky130_fd_sc_hd__a31o_1 c687 (.A1(net523),
    .A2(net812),
    .A3(clknet_1_1__leaf_net532),
    .B1(clknet_1_0__leaf_net742),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(clknet_1_1__leaf_net521),
    .A1(clknet_1_0__leaf_net436),
    .A2(net534),
    .A3(clknet_1_0__leaf_net538),
    .S0(clknet_1_0__leaf_net518),
    .S1(clknet_1_0__leaf_net535),
    .X(net541));
 sky130_fd_sc_hd__sedfxbp_1 c689 (.CLK(clknet_4_1_0_clk),
    .D(net918),
    .DE(clknet_1_1__leaf_net436),
    .SCD(net524),
    .SCE(net707),
    .Q(net542));
 sky130_fd_sc_hd__xnor2_4 c69 (.A(net840),
    .B(net807),
    .Y(net7));
 sky130_fd_sc_hd__sdfbbn_1 c690 (.CLK_N(clknet_4_0_0_clk),
    .D(clknet_1_0__leaf_net519),
    .RESET_B(clknet_1_0__leaf_net538),
    .SCD(net515),
    .SCE(net218),
    .SET_B(clknet_1_0__leaf_net742),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__a31o_1 c691 (.A1(net97),
    .A2(net427),
    .A3(net669),
    .B1(clknet_1_0__leaf_net742),
    .X(net545));
 sky130_fd_sc_hd__sdfbbn_1 c692 (.CLK_N(clknet_4_1_0_clk),
    .D(net332),
    .RESET_B(clknet_1_1__leaf_net529),
    .SCD(clknet_1_1__leaf_net519),
    .SCE(net908),
    .SET_B(net533),
    .Q(net547),
    .Q_N(net546));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(clknet_1_0__leaf_net537),
    .A1(net903),
    .A2(net543),
    .A3(clknet_1_0__leaf_net535),
    .S0(clknet_1_0__leaf_net521),
    .S1(clknet_1_0__leaf_net436),
    .X(net548));
 sky130_fd_sc_hd__a31o_1 c694 (.A1(net223),
    .A2(clknet_1_0__leaf_net538),
    .A3(net544),
    .B1(net546),
    .X(net549));
 sky130_fd_sc_hd__a31o_1 c695 (.A1(net547),
    .A2(clknet_1_0__leaf_net535),
    .A3(net669),
    .B1(clknet_1_0__leaf_net742),
    .X(net550));
 sky130_fd_sc_hd__a41o_1 c696 (.A1(clknet_1_1__leaf_net545),
    .A2(clknet_1_0__leaf_net521),
    .A3(net223),
    .A4(net427),
    .B1(net709),
    .X(net551));
 sky130_fd_sc_hd__sedfxtp_1 c697 (.CLK(clknet_4_0_0_clk),
    .D(net515),
    .DE(net218),
    .SCD(clknet_1_0__leaf_net548),
    .SCE(net523),
    .Q(net552));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(clknet_1_0__leaf_net408),
    .A2(clknet_1_0__leaf_net545),
    .A3(net552),
    .B1(clknet_1_0__leaf_net537),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_1__leaf_net551),
    .A1(net97),
    .A2(net523),
    .A3(clknet_1_1__leaf_net529),
    .S0(clknet_1_1__leaf_net550),
    .S1(net929),
    .X(net554));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net6),
    .B(net4),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net544),
    .A1(net413),
    .A2(net552),
    .A3(clknet_1_0__leaf_net553),
    .S0(clknet_1_0__leaf_net551),
    .S1(clknet_1_0__leaf_net742),
    .X(net555));
 sky130_fd_sc_hd__a41o_1 c701 (.A1(clknet_1_1__leaf_net540),
    .A2(clknet_1_0__leaf_net550),
    .A3(clknet_1_0__leaf_net545),
    .A4(clknet_1_1__leaf_net436),
    .B1(net530),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net555),
    .A1(net552),
    .A2(clknet_1_1__leaf_net556),
    .A3(net429),
    .S0(net918),
    .S1(clknet_1_0__leaf_net540),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net221),
    .A1(clknet_1_0__leaf_net556),
    .A2(clknet_1_0__leaf_net554),
    .A3(clknet_1_0__leaf_net550),
    .S0(clknet_1_0__leaf_net551),
    .S1(net743),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net413),
    .A1(net218),
    .A2(net842),
    .A3(clknet_1_1__leaf_net535),
    .S0(net923),
    .S1(clknet_1_1__leaf_net742),
    .X(net559));
 sky130_fd_sc_hd__sdfbbp_1 c705 (.CLK(clknet_4_3_0_clk),
    .D(net430),
    .RESET_B(net845),
    .SCD(clknet_1_0__leaf_net459),
    .SCE(net524),
    .SET_B(net837),
    .Q(net561),
    .Q_N(net560));
 sky130_fd_sc_hd__a41o_1 c706 (.A1(clknet_1_1__leaf_net554),
    .A2(net524),
    .A3(net238),
    .A4(net561),
    .B1(net530),
    .X(net562));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_0_0_clk),
    .D(net333),
    .RESET_B(net218),
    .SCD(net561),
    .SCE(net812),
    .SET_B(clknet_1_0__leaf_net742),
    .Q(net564),
    .Q_N(net563));
 sky130_fd_sc_hd__a41o_1 c708 (.A1(net837),
    .A2(net564),
    .A3(net560),
    .A4(clknet_1_0__leaf_net742),
    .B1(net745),
    .X(net565));
 sky130_fd_sc_hd__sdfbbn_1 c709 (.CLK_N(clknet_4_0_0_clk),
    .D(net524),
    .RESET_B(net794),
    .SCD(net534),
    .SCE(clknet_1_0__leaf_net548),
    .SET_B(net560),
    .Q(net566));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net825),
    .B(net842),
    .Y(net9));
 sky130_fd_sc_hd__sdfbbp_1 c710 (.CLK(clknet_4_2_0_clk),
    .D(net327),
    .RESET_B(clknet_1_1__leaf_net548),
    .SCD(net533),
    .SCE(net413),
    .SET_B(net729),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__sdfbbn_1 c711 (.CLK_N(clknet_4_2_0_clk),
    .D(clknet_1_1__leaf_net556),
    .RESET_B(net929),
    .SCD(net534),
    .SCE(net563),
    .SET_B(net561),
    .Q(net570),
    .Q_N(net569));
 sky130_fd_sc_hd__sdfbbn_1 c712 (.CLK_N(clknet_4_2_0_clk),
    .D(net968),
    .RESET_B(clknet_1_0__leaf_net548),
    .SCD(clknet_1_0__leaf_net449),
    .SCE(net561),
    .SET_B(net935),
    .Q(net571));
 sky130_fd_sc_hd__a41o_1 c713 (.A1(net542),
    .A2(net106),
    .A3(net533),
    .A4(net563),
    .B1(net937),
    .X(net572));
 sky130_fd_sc_hd__a41o_1 c714 (.A1(net561),
    .A2(net571),
    .A3(net903),
    .A4(net533),
    .B1(net77),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net573),
    .A1(net238),
    .A2(net799),
    .A3(net560),
    .S0(clknet_1_1__leaf_net742),
    .S1(net744),
    .X(net574));
 sky130_fd_sc_hd__sdfbbp_1 c716 (.CLK(clknet_4_0_0_clk),
    .D(net566),
    .RESET_B(net572),
    .SCD(clknet_1_0__leaf_net554),
    .SCE(net429),
    .SET_B(net935),
    .Q(net575));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(clknet_1_1__leaf_net553),
    .A1(net572),
    .A2(net573),
    .A3(net837),
    .S0(net935),
    .S1(net747),
    .X(net576));
 sky130_fd_sc_hd__sdfbbn_1 c718 (.CLK_N(clknet_4_0_0_clk),
    .D(net565),
    .RESET_B(net534),
    .SCD(net908),
    .SCE(net524),
    .SET_B(net923),
    .Q(net578),
    .Q_N(net577));
 sky130_fd_sc_hd__sdfbbn_1 c719 (.CLK_N(clknet_4_0_0_clk),
    .D(net908),
    .RESET_B(clknet_1_0__leaf_net556),
    .SCD(net560),
    .SCE(net745),
    .SET_B(net748),
    .Q(net579));
 sky130_fd_sc_hd__xnor2_4 c72 (.A(net823),
    .B(net936),
    .Y(net10));
 sky130_fd_sc_hd__a41o_1 c720 (.A1(net575),
    .A2(net572),
    .A3(net77),
    .A4(net238),
    .B1(net746),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net579),
    .A1(net580),
    .A2(net791),
    .A3(net218),
    .S0(net856),
    .S1(net935),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net578),
    .A1(net572),
    .A2(net567),
    .A3(net812),
    .S0(net837),
    .S1(net560),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net549),
    .A1(net570),
    .A2(net937),
    .A3(clknet_1_1__leaf_net548),
    .S0(net577),
    .S1(net935),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net218),
    .A1(clknet_1_0__leaf_net449),
    .A2(net569),
    .A3(net244),
    .S0(net561),
    .S1(net396),
    .X(net584));
 sky130_fd_sc_hd__sdfbbp_1 c725 (.CLK(clknet_4_2_0_clk),
    .D(clknet_1_1__leaf_net548),
    .RESET_B(net582),
    .SCD(net560),
    .SCE(net749),
    .SET_B(net960),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net582),
    .A1(net530),
    .A2(clknet_1_1__leaf_net535),
    .A3(net238),
    .S0(net710),
    .S1(net747),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net396),
    .A1(net932),
    .A2(net467),
    .A3(net546),
    .S0(net746),
    .S1(net750),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net547),
    .A1(net837),
    .A2(net430),
    .A3(clknet_1_0__leaf_net486),
    .S0(net79),
    .S1(net912),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net459),
    .A1(net908),
    .A2(net244),
    .A3(net733),
    .S0(clknet_1_1__leaf_net742),
    .S1(net746),
    .X(net590));
 sky130_fd_sc_hd__xnor2_4 c73 (.A(net847),
    .B(net2),
    .Y(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net106),
    .A1(net396),
    .A2(net908),
    .A3(clknet_1_1__leaf_net535),
    .S0(net712),
    .S1(net751),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net106),
    .A1(net932),
    .A2(net430),
    .A3(net915),
    .S0(net473),
    .S1(net913),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(clknet_1_0__leaf_net479),
    .A1(net588),
    .A2(net547),
    .A3(net468),
    .S0(net908),
    .S1(clknet_1_1__leaf_net535),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net530),
    .A1(clknet_1_0__leaf_net486),
    .A2(net923),
    .A3(clknet_1_1__leaf_net742),
    .S0(net747),
    .S1(net752),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net535),
    .A1(net250),
    .A2(net915),
    .A3(net923),
    .S0(clknet_1_1__leaf_net742),
    .S1(net746),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net250),
    .A1(net915),
    .A2(net932),
    .A3(net908),
    .S0(net730),
    .S1(clknet_1_1__leaf_net742),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net923),
    .A1(net596),
    .A2(net908),
    .A3(clknet_1_1__leaf_net591),
    .S0(net472),
    .S1(net746),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net908),
    .A1(net594),
    .A2(net905),
    .A3(net932),
    .S0(net915),
    .S1(net796),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net110),
    .A1(clknet_1_0__leaf_net597),
    .A2(net530),
    .A3(net788),
    .S1(net729),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(clknet_1_1__leaf_net459),
    .A1(net589),
    .A2(clknet_1_0__leaf_net597),
    .A3(net923),
    .S0(net546),
    .S1(net747),
    .X(net600));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net2),
    .B(net9),
    .Y(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net592),
    .A1(net590),
    .A2(net322),
    .A3(net923),
    .S0(net934),
    .S1(net746),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net592),
    .A1(net473),
    .A2(clknet_1_0__leaf_net597),
    .A3(net530),
    .S0(net747),
    .S1(net752),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(net876),
    .A1(clknet_1_0__leaf_net597),
    .A2(net672),
    .A3(net747),
    .S0(net753),
    .S1(net756),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_0__leaf_net591),
    .A1(net527),
    .A2(net430),
    .A3(net905),
    .S0(net754),
    .S1(net755),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net110),
    .A1(clknet_1_0__leaf_net597),
    .A2(net592),
    .A3(net795),
    .S0(net683),
    .S1(net757),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net601),
    .A1(net604),
    .A2(net530),
    .A3(net913),
    .S0(clknet_1_0__leaf_net597),
    .S1(net758),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net322),
    .A1(net595),
    .A2(net396),
    .A3(net585),
    .S0(net758),
    .S1(net759),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net587),
    .A1(net607),
    .A2(net918),
    .A3(clknet_1_1__leaf_net597),
    .S0(net758),
    .S1(net759),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net904),
    .A1(clknet_1_1__leaf_net597),
    .A2(net392),
    .A3(clknet_1_1__leaf_net474),
    .S0(net937),
    .S1(net708),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net238),
    .A1(net392),
    .A2(clknet_1_1__leaf_net538),
    .A3(net79),
    .S0(clknet_1_1__leaf_net597),
    .S1(clknet_1_0__leaf_net761),
    .X(net610));
 sky130_fd_sc_hd__xnor2_4 c75 (.A(net11),
    .B(net10),
    .Y(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_1__leaf_net538),
    .A1(net77),
    .A2(clknet_1_1__leaf_net486),
    .A3(net904),
    .S0(net935),
    .S1(clknet_1_0__leaf_net741),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net934),
    .A1(clknet_1_1__leaf_net538),
    .A2(net392),
    .A3(clknet_1_1__leaf_net741),
    .S0(clknet_1_1__leaf_net760),
    .S1(clknet_1_1__leaf_net761),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_1__leaf_net474),
    .A1(clknet_1_1__leaf_net511),
    .A2(net392),
    .A3(net660),
    .S0(net708),
    .S1(clknet_1_0__leaf_net760),
    .X(net613));
 sky130_fd_sc_hd__mux4_2 c753 (.A0(net568),
    .A1(net586),
    .A2(clknet_1_0__leaf_net511),
    .A3(net467),
    .S0(net812),
    .S1(clknet_1_0__leaf_net760),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net905),
    .A1(net530),
    .A2(net913),
    .A3(clknet_1_1__leaf_net474),
    .S0(net392),
    .S1(clknet_1_1__leaf_net762),
    .X(net615));
 sky130_fd_sc_hd__mux4_2 c755 (.A0(net473),
    .A1(net614),
    .A2(net856),
    .A3(net934),
    .S0(net708),
    .S1(clknet_1_0__leaf_net762),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net913),
    .A1(net611),
    .A2(net392),
    .A3(net470),
    .S0(net244),
    .S1(net812),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net934),
    .A1(net904),
    .A2(net392),
    .A3(net731),
    .S0(net767),
    .S1(net768),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net876),
    .A1(clknet_1_1__leaf_net597),
    .A2(net79),
    .A3(net671),
    .S0(net767),
    .S1(net769),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(clknet_1_1__leaf_net486),
    .A1(net470),
    .A2(net904),
    .A3(net731),
    .S0(net766),
    .S1(net769),
    .X(net620));
 sky130_fd_sc_hd__mux4_2 c76 (.A0(net807),
    .A1(net798),
    .A2(net839),
    .A3(net8),
    .S0(net12),
    .S1(net832),
    .X(net14));
 sky130_fd_sc_hd__mux4_2 c760 (.A0(net238),
    .A1(clknet_1_0__leaf_net511),
    .A2(net708),
    .A3(net764),
    .S0(net766),
    .S1(net770),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net530),
    .A1(net933),
    .A2(net913),
    .A3(clknet_1_0__leaf_net741),
    .S0(net768),
    .S1(net770),
    .X(net622));
 sky130_fd_sc_hd__mux4_2 c762 (.A0(net468),
    .A1(net621),
    .A2(clknet_1_1__leaf_net622),
    .A3(net933),
    .S0(clknet_1_1__leaf_net741),
    .S1(net765),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(clknet_1_0__leaf_net620),
    .A1(net933),
    .A2(net110),
    .A3(net530),
    .S0(net677),
    .S1(net771),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(clknet_1_0__leaf_net622),
    .A1(clknet_1_1__leaf_net620),
    .A2(net913),
    .A3(net697),
    .S0(clknet_1_0__leaf_net741),
    .S1(net763),
    .X(net625));
 sky130_fd_sc_hd__xnor2_4 c77 (.A(net14),
    .B(net5),
    .Y(net15));
 sky130_fd_sc_hd__mux4_2 c78 (.A0(net835),
    .A1(net841),
    .A2(net844),
    .A3(net12),
    .S0(net15),
    .S1(net14),
    .X(net16));
 sky130_fd_sc_hd__xnor2_4 c79 (.A(net936),
    .B(net930),
    .Y(net864));
 sky130_fd_sc_hd__xnor2_4 c80 (.A(net826),
    .B(net7),
    .Y(net17));
 sky130_fd_sc_hd__xnor2_4 c81 (.A(net17),
    .B(net16),
    .Y(net18));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net10),
    .A1(net7),
    .A2(net936),
    .A3(net922),
    .S0(net12),
    .S1(net15),
    .X(net19));
 sky130_fd_sc_hd__xnor2_2 c83 (.A(net17),
    .B(net832),
    .Y(net20));
 sky130_fd_sc_hd__xnor2_2 c84 (.A(net18),
    .B(net4),
    .Y(net21));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net8),
    .A1(net9),
    .A2(net21),
    .A3(net12),
    .S0(net805),
    .S1(net15),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net21),
    .A1(net11),
    .A2(net18),
    .A3(net19),
    .S0(net13),
    .S1(net22),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net830),
    .A1(net23),
    .A2(net22),
    .A3(net936),
    .S0(net804),
    .S1(net922),
    .X(net24));
 sky130_fd_sc_hd__xnor2_4 c88 (.A(net804),
    .B(net847),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_1 c89 (.A(net10),
    .B(net16),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net812),
    .B(net8),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_4 c91 (.A(net827),
    .B(net13),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_2 c92 (.A(net27),
    .B(net20),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net841),
    .B(net27),
    .Y(net30));
 sky130_fd_sc_hd__a41o_1 c94 (.A1(net22),
    .A2(net28),
    .A3(net29),
    .A4(net20),
    .B1(net30),
    .X(net31));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net30),
    .B(net864),
    .Y(net32));
 sky130_fd_sc_hd__a21bo_1 c96 (.A1(net13),
    .A2(net14),
    .B1_N(net27),
    .X(net33));
 sky130_fd_sc_hd__a21bo_1 c97 (.A1(net29),
    .A2(net33),
    .B1_N(net30),
    .X(net34));
 sky130_fd_sc_hd__mux4_2 c98 (.A0(net34),
    .A1(net834),
    .A2(net33),
    .A3(net930),
    .S0(net32),
    .S1(net28),
    .X(net35));
 sky130_fd_sc_hd__a21bo_4 c99 (.A1(net31),
    .A2(net35),
    .B1_N(net28),
    .X(net36));
 sky130_fd_sc_hd__a31o_1 merge765 (.A1(clknet_1_1__leaf_net518),
    .A2(net524),
    .A3(clknet_1_1__leaf_net528),
    .B1(clknet_1_0__leaf_net724),
    .X(net626));
 sky130_fd_sc_hd__a31o_1 merge766 (.A1(net233),
    .A2(net210),
    .A3(net232),
    .B1(net237),
    .X(net627));
 sky130_fd_sc_hd__a41o_1 merge767 (.A1(net18),
    .A2(net917),
    .A3(net124),
    .A4(net112),
    .B1(net833),
    .X(net628));
 sky130_fd_sc_hd__a31o_1 merge768 (.A1(net350),
    .A2(clknet_1_1__leaf_net431),
    .A3(net831),
    .B1(clknet_1_0__leaf_net416),
    .X(net629));
 sky130_fd_sc_hd__a41o_1 merge769 (.A1(net319),
    .A2(net312),
    .A3(net323),
    .A4(net318),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net161),
    .A1(net941),
    .A2(net839),
    .A3(net211),
    .S0(clknet_1_1__leaf_net269),
    .S1(net905),
    .X(net631));
 sky130_fd_sc_hd__mux4_2 merge771 (.A0(net157),
    .A1(net161),
    .A2(net132),
    .A3(net158),
    .S0(net904),
    .X(net662));
 sky130_fd_sc_hd__a41o_1 merge772 (.A1(net316),
    .A2(net337),
    .A3(net312),
    .A4(net293),
    .B1(net333),
    .X(net633));
 sky130_fd_sc_hd__a41o_1 merge773 (.A1(clknet_1_0__leaf_net406),
    .A2(clknet_1_0__leaf_net411),
    .A3(clknet_1_0__leaf_net412),
    .A4(net929),
    .B1(net398),
    .X(net634));
 sky130_fd_sc_hd__a41o_1 merge774 (.A1(net199),
    .A2(net216),
    .A3(net211),
    .A4(net219),
    .B1(net964),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net292),
    .A1(net266),
    .A2(net138),
    .A3(net122),
    .S0(net354),
    .S1(net219),
    .X(net636));
 sky130_fd_sc_hd__a31o_1 merge776 (.A1(clknet_1_1__leaf_net412),
    .A2(clknet_1_1__leaf_net408),
    .A3(clknet_1_0__leaf_net421),
    .B1(net424),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net789),
    .A1(net234),
    .A2(net250),
    .A3(net252),
    .S0(net138),
    .S1(net122),
    .X(net638));
 sky130_fd_sc_hd__a31o_1 merge778 (.A1(net55),
    .A2(net54),
    .A3(net137),
    .B1(net168),
    .X(net639));
 sky130_fd_sc_hd__a41o_1 merge779 (.A1(net101),
    .A2(net114),
    .A3(net360),
    .A4(net715),
    .B1(net716),
    .X(net640));
 sky130_fd_sc_hd__a41o_1 merge780 (.A1(net404),
    .A2(net424),
    .A3(net426),
    .A4(clknet_1_0__leaf_net428),
    .B1(net417),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net424),
    .A1(clknet_1_1__leaf_net531),
    .A2(clknet_1_1__leaf_net518),
    .A3(net522),
    .S0(clknet_1_0__leaf_net706),
    .S1(net725),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(clknet_1_1__leaf_net423),
    .A1(net903),
    .A2(net445),
    .A3(net228),
    .S0(net233),
    .S1(net232),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net354),
    .A1(net872),
    .A2(net360),
    .A3(net666),
    .S0(net696),
    .S1(net715),
    .X(net644));
 sky130_fd_sc_hd__sdfbbn_1 merge784 (.CLK_N(clknet_4_12_0_clk),
    .D(net163),
    .RESET_B(net145),
    .SCD(net274),
    .SCE(net162),
    .SET_B(net135),
    .Q(net646),
    .Q_N(net645));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net66),
    .A1(net229),
    .A2(net218),
    .A3(net973),
    .S0(net234),
    .S1(net959),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net177),
    .A1(net128),
    .A2(net900),
    .A3(net282),
    .S0(net850),
    .S1(net670),
    .X(net648));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net281),
    .A1(net282),
    .A2(net946),
    .A3(net258),
    .S0(net110),
    .S1(net884),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net403),
    .A1(net417),
    .A2(net811),
    .A3(net424),
    .S0(net309),
    .S1(net297),
    .X(net650));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(clknet_1_0__leaf_net419),
    .A1(clknet_1_1__leaf_net412),
    .A2(net921),
    .A3(clknet_1_0__leaf_net457),
    .S0(net935),
    .S1(net851),
    .X(net651));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net357),
    .A1(net360),
    .A2(net325),
    .A3(net234),
    .S0(net865),
    .S1(net947),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net439),
    .A1(clknet_1_1__leaf_net416),
    .A2(net333),
    .A3(net229),
    .S0(net238),
    .S1(net241),
    .X(net653));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net204),
    .A1(net211),
    .A2(net112),
    .A3(net283),
    .S0(net128),
    .S1(net680),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net250),
    .A1(net229),
    .A2(net234),
    .A3(clknet_1_1__leaf_net416),
    .S0(net236),
    .S1(net912),
    .X(net655));
 sky130_fd_sc_hd__dfrbp_1 merge794 (.CLK(clknet_4_15_0_clk),
    .D(net56),
    .Q(net58),
    .Q_N(net656));
 sky130_fd_sc_hd__dfrbp_1 merge795 (.CLK(clknet_4_12_0_clk),
    .D(net355),
    .RESET_B(net370),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dfrtn_1 merge796 (.CLK_N(clknet_4_10_0_clk),
    .D(net625),
    .RESET_B(net612),
    .Q(net660));
 sky130_fd_sc_hd__dfrtp_1 merge797 (.CLK(clknet_4_9_0_clk),
    .D(net490),
    .RESET_B(net501),
    .Q(net661));
 sky130_fd_sc_hd__dfrtp_4 merge798 (.CLK(clknet_4_15_0_clk),
    .RESET_B(net164),
    .Q(net662));
 sky130_fd_sc_hd__dfrtp_4 merge799 (.CLK(clknet_4_1_0_clk),
    .D(net634),
    .RESET_B(net414),
    .Q(net663));
 sky130_fd_sc_hd__dfsbp_1 merge800 (.CLK(clknet_4_1_0_clk),
    .D(net525),
    .SET_B(net626),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfsbp_1 merge801 (.CLK(clknet_4_6_0_clk),
    .D(net351),
    .Q(net352),
    .Q_N(net666));
 sky130_fd_sc_hd__dfstp_1 merge802 (.CLK(clknet_4_4_0_clk),
    .SET_B(net321),
    .Q(net630));
 sky130_fd_sc_hd__dfstp_1 merge803 (.CLK(clknet_4_1_0_clk),
    .D(net536),
    .SET_B(net541),
    .Q(net669));
 sky130_fd_sc_hd__dfstp_1 merge804 (.CLK(clknet_4_15_0_clk),
    .D(net275),
    .SET_B(net273),
    .Q(net670));
 sky130_fd_sc_hd__dlrbn_1 merge805 (.D(net559),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net562),
    .Q(net672),
    .Q_N(net671));
 sky130_fd_sc_hd__dlrbn_1 merge806 (.D(net179),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net180),
    .Q(net902),
    .Q_N(net673));
 sky130_fd_sc_hd__dlrbp_1 merge807 (.D(net268),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net255),
    .Q(net675),
    .Q_N(net674));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net144),
    .B(net140),
    .Y(net676));
 sky130_fd_sc_hd__dlrbp_1 merge809 (.D(net483),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net487),
    .Q(net678),
    .Q_N(net677));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net213),
    .B(net226),
    .Y(net679));
 sky130_fd_sc_hd__dlrtn_1 merge811 (.D(net242),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net627),
    .Q(net680));
 sky130_fd_sc_hd__xnor2_1 merge812 (.A(net441),
    .B(net452),
    .Y(net681));
 sky130_fd_sc_hd__dlrtn_1 merge813 (.D(net637),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net641),
    .Q(net682));
 sky130_fd_sc_hd__dlrtn_1 merge814 (.D(net373),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net379),
    .Q(net866));
 sky130_fd_sc_hd__dlrtp_1 merge815 (.D(net598),
    .GATE(clknet_4_8_0_clk),
    .Q(net599));
 sky130_fd_sc_hd__dlrtp_1 merge816 (.GATE(clknet_4_15_0_clk),
    .RESET_B(net289),
    .Q(net290));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net227),
    .B(net263),
    .Y(net684));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net488),
    .B(net624),
    .Y(net685));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net640),
    .B(net628),
    .Y(net686));
 sky130_fd_sc_hd__dlrtp_2 merge820 (.D(net676),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net686),
    .Q(net687));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net635),
    .B(net679),
    .Y(net688));
 sky130_fd_sc_hd__edfxbp_1 merge822 (.CLK(clknet_4_6_0_clk),
    .D(net633),
    .DE(net353),
    .Q(net690),
    .Q_N(net689));
 sky130_fd_sc_hd__edfxtp_1 merge823 (.CLK(clknet_4_14_0_clk),
    .D(net383),
    .DE(net184),
    .Q(net691));
 sky130_fd_sc_hd__sdlclkp_1 merge824 (.CLK(clknet_4_15_0_clk),
    .GATE(net183),
    .SCE(net639),
    .GCLK(net898));
 sky130_fd_sc_hd__sdlclkp_2 merge825 (.CLK(clknet_4_12_0_clk),
    .GATE(net652),
    .SCE(net644),
    .GCLK(net692));
 sky130_fd_sc_hd__sdlclkp_4 merge826 (.CLK(clknet_4_3_0_clk),
    .GATE(net681),
    .SCE(net642),
    .GCLK(net693));
 sky130_fd_sc_hd__dfrbp_1 merge827 (.CLK(clknet_4_14_0_clk),
    .D(net276),
    .RESET_B(net286),
    .Q(net694),
    .Q_N(net863));
 sky130_fd_sc_hd__dfrbp_1 merge828 (.CLK(clknet_4_13_0_clk),
    .D(net270),
    .RESET_B(net647),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__dfrtn_1 merge829 (.CLK_N(clknet_4_9_0_clk),
    .D(net685),
    .RESET_B(net629),
    .Q(net697));
 sky130_fd_sc_hd__dfrtp_4 merge830 (.CLK(clknet_4_5_0_clk),
    .D(net215),
    .RESET_B(net684),
    .Q(net698));
 sky130_fd_sc_hd__dfrtp_4 merge831 (.CLK(clknet_4_5_0_clk),
    .D(net205),
    .RESET_B(net688),
    .Q(net699));
 sky130_fd_sc_hd__dfxbp_1 s832 (.CLK(clknet_4_15_0_clk),
    .D(net57),
    .Q(net897),
    .Q_N(net700));
 sky130_fd_sc_hd__dfxbp_1 s833 (.CLK(clknet_4_7_0_clk),
    .D(net139),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__dfxtp_2 s834 (.CLK(clknet_4_5_0_clk),
    .D(net212),
    .Q(net703));
 sky130_fd_sc_hd__dfxtp_4 s835 (.CLK(clknet_4_5_0_clk),
    .D(net224),
    .Q(net704));
 sky130_fd_sc_hd__dfxtp_1 s836 (.CLK(clknet_4_13_0_clk),
    .D(net264),
    .Q(net705));
 sky130_fd_sc_hd__dlclkp_1 s837 (.CLK(clknet_4_14_0_clk),
    .GATE(net287),
    .GCLK(net874));
 sky130_fd_sc_hd__dlclkp_2 s838 (.CLK(clknet_4_15_0_clk),
    .GATE(net288),
    .GCLK(net854));
 sky130_fd_sc_hd__dlclkp_4 s839 (.CLK(clknet_4_4_0_clk),
    .GATE(net324),
    .GCLK(net706));
 sky130_fd_sc_hd__dlxbn_2 s840 (.D(net326),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net708),
    .Q_N(net707));
 sky130_fd_sc_hd__dlxbn_2 s841 (.D(net329),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dlxbp_1 s842 (.D(net331),
    .GATE(clknet_4_4_0_clk),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dlxtn_1 s843 (.D(net346),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net713));
 sky130_fd_sc_hd__dlxtn_1 s844 (.D(net348),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net714));
 sky130_fd_sc_hd__dlxtn_2 s845 (.D(net349),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net715));
 sky130_fd_sc_hd__dlxtp_1 s846 (.D(net363),
    .GATE(clknet_4_13_0_clk),
    .Q(net716));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s847 (.D(net369),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net717));
 sky130_fd_sc_hd__dfxbp_1 s848 (.CLK(clknet_4_14_0_clk),
    .D(net381),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dfxbp_1 s849 (.CLK(clknet_4_14_0_clk),
    .D(net382),
    .Q(net867));
 sky130_fd_sc_hd__dfxtp_1 s850 (.CLK(clknet_4_9_0_clk),
    .D(net384),
    .Q(net720));
 sky130_fd_sc_hd__dfxtp_2 s851 (.CLK(clknet_4_14_0_clk),
    .D(net386),
    .Q(net721));
 sky130_fd_sc_hd__dfxtp_1 s852 (.CLK(clknet_4_14_0_clk),
    .D(net390),
    .Q(net722));
 sky130_fd_sc_hd__dlclkp_1 s853 (.CLK(clknet_4_14_0_clk),
    .GATE(net391),
    .GCLK(net723));
 sky130_fd_sc_hd__dlclkp_2 s854 (.CLK(clknet_4_11_0_clk),
    .GATE(net393),
    .GCLK(net883));
 sky130_fd_sc_hd__dlclkp_4 s855 (.CLK(clknet_4_4_0_clk),
    .GATE(net405),
    .GCLK(net724));
 sky130_fd_sc_hd__dlxbn_1 s856 (.D(net432),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__dlxbn_1 s857 (.D(net434),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dlxbp_1 s858 (.D(net438),
    .GATE(clknet_4_1_0_clk),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlxtn_1 s859 (.D(net454),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net731));
 sky130_fd_sc_hd__dlxtn_1 s860 (.D(net456),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net851));
 sky130_fd_sc_hd__dlxtn_1 s861 (.D(net458),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net732));
 sky130_fd_sc_hd__dlxtp_1 s862 (.D(net478),
    .GATE(clknet_4_3_0_clk),
    .Q(net880));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s863 (.D(net482),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net733));
 sky130_fd_sc_hd__dfxbp_1 s864 (.CLK(clknet_4_9_0_clk),
    .D(net484),
    .Q(net735),
    .Q_N(net734));
 sky130_fd_sc_hd__dfxbp_2 s865 (.CLK(clknet_4_11_0_clk),
    .D(net499),
    .Q(net870),
    .Q_N(net736));
 sky130_fd_sc_hd__dfxtp_1 s866 (.CLK(clknet_4_11_0_clk),
    .D(net500),
    .Q(net737));
 sky130_fd_sc_hd__dfxtp_1 s867 (.CLK(clknet_4_11_0_clk),
    .D(net505),
    .Q(net738));
 sky130_fd_sc_hd__dfxtp_1 s868 (.CLK(clknet_4_11_0_clk),
    .D(net507),
    .Q(net739));
 sky130_fd_sc_hd__dlclkp_1 s869 (.CLK(clknet_4_11_0_clk),
    .GATE(net508),
    .GCLK(net740));
 sky130_fd_sc_hd__dlclkp_2 s870 (.CLK(clknet_4_10_0_clk),
    .GATE(net510),
    .GCLK(net741));
 sky130_fd_sc_hd__dlclkp_4 s871 (.CLK(clknet_4_0_0_clk),
    .GATE(net539),
    .GCLK(net742));
 sky130_fd_sc_hd__dlxbn_1 s872 (.D(net557),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxbn_1 s873 (.D(net558),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dlxbp_1 s874 (.D(net574),
    .GATE(clknet_4_2_0_clk),
    .Q(net747),
    .Q_N(net746));
 sky130_fd_sc_hd__dlxtn_1 s875 (.D(net576),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net748));
 sky130_fd_sc_hd__dlxtn_1 s876 (.D(net581),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__dlxtn_1 s877 (.D(net583),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net750));
 sky130_fd_sc_hd__dlxtp_1 s878 (.D(net584),
    .GATE(clknet_4_3_0_clk),
    .Q(net751));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s879 (.D(net593),
    .SLEEP_B(clknet_4_2_0_clk),
    .Q(net752));
 sky130_fd_sc_hd__dfxbp_1 s880 (.CLK(clknet_4_2_0_clk),
    .D(net600),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dfxbp_1 s881 (.CLK(clknet_4_2_0_clk),
    .D(net602),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__dfxtp_1 s882 (.CLK(clknet_4_8_0_clk),
    .D(net603),
    .Q(net757));
 sky130_fd_sc_hd__dfxtp_1 s883 (.CLK(clknet_4_8_0_clk),
    .D(net605),
    .Q(net758));
 sky130_fd_sc_hd__dfxtp_1 s884 (.CLK(clknet_4_8_0_clk),
    .D(net606),
    .Q(net759));
 sky130_fd_sc_hd__dlclkp_1 s885 (.CLK(clknet_4_8_0_clk),
    .GATE(net608),
    .GCLK(net760));
 sky130_fd_sc_hd__dlclkp_2 s886 (.CLK(clknet_4_10_0_clk),
    .GATE(net609),
    .GCLK(net761));
 sky130_fd_sc_hd__dlclkp_4 s887 (.CLK(clknet_4_8_0_clk),
    .GATE(net610),
    .GCLK(net762));
 sky130_fd_sc_hd__dlxbn_1 s888 (.D(net613),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxbn_1 s889 (.D(net615),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__dlxbp_1 s890 (.D(net616),
    .GATE(clknet_4_8_0_clk),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__dlxtn_1 s891 (.D(net617),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dlxtn_1 s892 (.D(net618),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net769));
 sky130_fd_sc_hd__dlxtn_1 s893 (.D(net619),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net770));
 sky130_fd_sc_hd__dlxtp_1 s894 (.D(net623),
    .GATE(clknet_4_10_0_clk),
    .Q(net771));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s895 (.D(net631),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net772));
 sky130_fd_sc_hd__dfxbp_1 s896 (.CLK(clknet_4_12_0_clk),
    .D(net636),
    .Q(net774),
    .Q_N(net773));
 sky130_fd_sc_hd__dfxbp_1 s897 (.CLK(clknet_4_13_0_clk),
    .D(net638),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__dfxtp_1 s898 (.CLK(clknet_4_5_0_clk),
    .D(net643),
    .Q(net777));
 sky130_fd_sc_hd__dfxtp_1 s899 (.CLK(clknet_4_15_0_clk),
    .D(net648),
    .Q(net778));
 sky130_fd_sc_hd__dfxtp_1 s900 (.CLK(clknet_4_15_0_clk),
    .D(net649),
    .Q(net779));
 sky130_fd_sc_hd__dlclkp_1 s901 (.CLK(clknet_4_4_0_clk),
    .GATE(net650),
    .GCLK(net780));
 sky130_fd_sc_hd__dlclkp_2 s902 (.CLK(clknet_4_1_0_clk),
    .GATE(net651),
    .GCLK(net781));
 sky130_fd_sc_hd__dlclkp_4 s903 (.CLK(clknet_4_7_0_clk),
    .GATE(net653),
    .GCLK(net782));
 sky130_fd_sc_hd__dlxbn_1 s904 (.D(net654),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__dlxbn_1 s905 (.D(net655),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net787));
 sky130_fd_sc_hd__buf_4 input3 (.A(in10),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net790));
 sky130_fd_sc_hd__buf_2 input6 (.A(in13),
    .X(net791));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net793));
 sky130_fd_sc_hd__buf_4 input9 (.A(in16),
    .X(net794));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net795));
 sky130_fd_sc_hd__buf_4 input11 (.A(in18),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net797));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net798));
 sky130_fd_sc_hd__buf_4 input14 (.A(in20),
    .X(net799));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net800));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net801));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_8 input19 (.A(in25),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in28),
    .X(net807));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net808));
 sky130_fd_sc_hd__buf_2 input24 (.A(in3),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(in31),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_8 input27 (.A(in32),
    .X(net812));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net816));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net819));
 sky130_fd_sc_hd__buf_2 input35 (.A(in4),
    .X(net820));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in43),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in44),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net827));
 sky130_fd_sc_hd__buf_2 input43 (.A(in47),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net830));
 sky130_fd_sc_hd__buf_2 input46 (.A(in5),
    .X(net831));
 sky130_fd_sc_hd__buf_4 input47 (.A(in50),
    .X(net832));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net833));
 sky130_fd_sc_hd__buf_4 input49 (.A(in52),
    .X(net834));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net835));
 sky130_fd_sc_hd__buf_8 input51 (.A(in54),
    .X(net836));
 sky130_fd_sc_hd__buf_4 input52 (.A(in55),
    .X(net837));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(in57),
    .X(net839));
 sky130_fd_sc_hd__buf_4 input55 (.A(in58),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(in6),
    .X(net842));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net844));
 sky130_fd_sc_hd__buf_4 input60 (.A(in7),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in8),
    .X(net846));
 sky130_fd_sc_hd__buf_4 input62 (.A(in9),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net848),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net849),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net850),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net851),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net852),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net853),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(clknet_1_1__leaf_net854),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net855),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net856),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output72 (.A(net934),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net858),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net859),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(clknet_1_1__leaf_net860),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(clknet_1_1__leaf_net861),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(clknet_1_1__leaf_net862),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output78 (.A(net863),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net864),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output80 (.A(net865),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output81 (.A(net866),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output82 (.A(net867),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net868),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output84 (.A(net920),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output85 (.A(net870),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net871),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net872),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(clknet_1_1__leaf_net873),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(clknet_1_1__leaf_net874),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net875),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output91 (.A(net876),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net877),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net878),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net879),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output95 (.A(net880),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net881),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net882),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net883),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net884),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net885),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net886),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net952),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net888),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output104 (.A(net889),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net890),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output106 (.A(net891),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(clknet_1_1__leaf_net892),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net893),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_1__leaf_net894),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net895),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net896),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net897),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(clknet_1_1__leaf_net898),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net899),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output115 (.A(net978),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output116 (.A(net901),
    .X(out8));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net902),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(net311),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net159),
    .X(net904));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net135),
    .X(net905));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net152),
    .X(net906));
 sky130_fd_sc_hd__buf_6 fanout122 (.A(net900),
    .X(net907));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net527),
    .X(net908));
 sky130_fd_sc_hd__buf_4 max_cap124 (.A(net848),
    .X(net909));
 sky130_fd_sc_hd__buf_4 max_cap125 (.A(net105),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net914),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net345),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net292),
    .X(net915));
 sky130_fd_sc_hd__buf_2 fanout131 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net85),
    .X(net918));
 sky130_fd_sc_hd__buf_4 max_cap134 (.A(net291),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net869),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net191),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net864),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net187),
    .X(net924));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net187),
    .X(net928));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(net75),
    .X(net929));
 sky130_fd_sc_hd__buf_4 max_cap145 (.A(net8),
    .X(net930));
 sky130_fd_sc_hd__buf_4 wire146 (.A(net67),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net934),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net857),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net731),
    .X(net935));
 sky130_fd_sc_hd__buf_4 max_cap151 (.A(net9),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net833),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net782 (.A(net782),
    .X(clknet_0_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net782 (.A(clknet_0_net782),
    .X(clknet_1_0__leaf_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net782 (.A(clknet_0_net782),
    .X(clknet_1_1__leaf_net782));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net449 (.A(net449),
    .X(clknet_0_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_0__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net449 (.A(clknet_0_net449),
    .X(clknet_1_1__leaf_net449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net243 (.A(net243),
    .X(clknet_0_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_0__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_1__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net257 (.A(net257),
    .X(clknet_0_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_0__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_1__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net262 (.A(net262),
    .X(clknet_0_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_0__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_1__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net269 (.A(net269),
    .X(clknet_0_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_0__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net269 (.A(clknet_0_net269),
    .X(clknet_1_1__leaf_net269));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net854 (.A(net854),
    .X(clknet_0_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_0__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net854 (.A(clknet_0_net854),
    .X(clknet_1_1__leaf_net854));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net894 (.A(net894),
    .X(clknet_0_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_0__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net894 (.A(clknet_0_net894),
    .X(clknet_1_1__leaf_net894));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net874 (.A(net874),
    .X(clknet_0_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_0__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net874 (.A(clknet_0_net874),
    .X(clknet_1_1__leaf_net874));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net265 (.A(net265),
    .X(clknet_0_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_0__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_1__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net781 (.A(net781),
    .X(clknet_0_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net781 (.A(clknet_0_net781),
    .X(clknet_1_0__leaf_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net781 (.A(clknet_0_net781),
    .X(clknet_1_1__leaf_net781));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net423 (.A(net423),
    .X(clknet_0_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_0__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net423 (.A(clknet_0_net423),
    .X(clknet_1_1__leaf_net423));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net537 (.A(net537),
    .X(clknet_0_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_0__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net537 (.A(clknet_0_net537),
    .X(clknet_1_1__leaf_net537));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net548 (.A(net548),
    .X(clknet_0_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_0__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_1__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net538 (.A(net538),
    .X(clknet_0_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_0__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_1__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net762 (.A(net762),
    .X(clknet_0_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net762 (.A(clknet_0_net762),
    .X(clknet_1_0__leaf_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net762 (.A(clknet_0_net762),
    .X(clknet_1_1__leaf_net762));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net433 (.A(net433),
    .X(clknet_0_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_0__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net433 (.A(clknet_0_net433),
    .X(clknet_1_1__leaf_net433));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net474 (.A(net474),
    .X(clknet_0_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_0__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net474 (.A(clknet_0_net474),
    .X(clknet_1_1__leaf_net474));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net761 (.A(net761),
    .X(clknet_0_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_0__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net761 (.A(clknet_0_net761),
    .X(clknet_1_1__leaf_net761));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net428 (.A(net428),
    .X(clknet_0_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_0__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_1__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net780 (.A(net780),
    .X(clknet_0_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_0__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net780 (.A(clknet_0_net780),
    .X(clknet_1_1__leaf_net780));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net431 (.A(net431),
    .X(clknet_0_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_0__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net431 (.A(clknet_0_net431),
    .X(clknet_1_1__leaf_net431));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net425 (.A(net425),
    .X(clknet_0_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_0__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net425 (.A(clknet_0_net425),
    .X(clknet_1_1__leaf_net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net760 (.A(net760),
    .X(clknet_0_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_1__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net550 (.A(net550),
    .X(clknet_0_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_0__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net550 (.A(clknet_0_net550),
    .X(clknet_1_1__leaf_net550));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net545 (.A(net545),
    .X(clknet_0_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_0__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_1__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net551 (.A(net551),
    .X(clknet_0_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_0__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_1__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net741 (.A(net741),
    .X(clknet_0_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_0__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_1__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net724 (.A(net724),
    .X(clknet_0_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_0__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_1__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net521 (.A(net521),
    .X(clknet_0_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_0__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net521 (.A(clknet_0_net521),
    .X(clknet_1_1__leaf_net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net520 (.A(net520),
    .X(clknet_0_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_0__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net520 (.A(clknet_0_net520),
    .X(clknet_1_1__leaf_net520));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net528 (.A(net528),
    .X(clknet_0_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net518 (.A(net518),
    .X(clknet_0_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_0__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net518 (.A(clknet_0_net518),
    .X(clknet_1_1__leaf_net518));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net513 (.A(net513),
    .X(clknet_0_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_0__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net513 (.A(clknet_0_net513),
    .X(clknet_1_1__leaf_net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net529 (.A(net529),
    .X(clknet_0_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net535 (.A(net535),
    .X(clknet_0_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_0__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net535 (.A(clknet_0_net535),
    .X(clknet_1_1__leaf_net535));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net591 (.A(net591),
    .X(clknet_0_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_0__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_1__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net531 (.A(net531),
    .X(clknet_0_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_0__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net531 (.A(clknet_0_net531),
    .X(clknet_1_1__leaf_net531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net519 (.A(net519),
    .X(clknet_0_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_0__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net519 (.A(clknet_0_net519),
    .X(clknet_1_1__leaf_net519));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net408 (.A(net408),
    .X(clknet_0_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_0__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net526 (.A(net526),
    .X(clknet_0_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_0__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net526 (.A(clknet_0_net526),
    .X(clknet_1_1__leaf_net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net406 (.A(net406),
    .X(clknet_0_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_0__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net406 (.A(clknet_0_net406),
    .X(clknet_1_1__leaf_net406));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net486 (.A(net486),
    .X(clknet_0_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_0__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net486 (.A(clknet_0_net486),
    .X(clknet_1_1__leaf_net486));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net620 (.A(net620),
    .X(clknet_0_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net620 (.A(clknet_0_net620),
    .X(clknet_1_0__leaf_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net620 (.A(clknet_0_net620),
    .X(clknet_1_1__leaf_net620));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net416 (.A(net416),
    .X(clknet_0_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_0__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_1__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net394 (.A(net394),
    .X(clknet_0_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_0__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net394 (.A(clknet_0_net394),
    .X(clknet_1_1__leaf_net394));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net706 (.A(net706),
    .X(clknet_0_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net419 (.A(net419),
    .X(clknet_0_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_0__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_1__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net692 (.A(net692),
    .X(clknet_0_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_0__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net692 (.A(clknet_0_net692),
    .X(clknet_1_1__leaf_net692));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net361 (.A(net361),
    .X(clknet_0_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_0__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net361 (.A(clknet_0_net361),
    .X(clknet_1_1__leaf_net361));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net362 (.A(net362),
    .X(clknet_0_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_0__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net362 (.A(clknet_0_net362),
    .X(clknet_1_1__leaf_net362));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net371 (.A(net371),
    .X(clknet_0_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_0__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net371 (.A(clknet_0_net371),
    .X(clknet_1_1__leaf_net371));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net860 (.A(net860),
    .X(clknet_0_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net860 (.A(clknet_0_net860),
    .X(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net862 (.A(net862),
    .X(clknet_0_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_0__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net862 (.A(clknet_0_net862),
    .X(clknet_1_1__leaf_net862));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net377 (.A(net377),
    .X(clknet_0_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_0__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net377 (.A(clknet_0_net377),
    .X(clknet_1_1__leaf_net377));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net861 (.A(net861),
    .X(clknet_0_net861));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net861 (.A(clknet_0_net861),
    .X(clknet_1_0__leaf_net861));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net861 (.A(clknet_0_net861),
    .X(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net364 (.A(net364),
    .X(clknet_0_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_0__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net364 (.A(clknet_0_net364),
    .X(clknet_1_1__leaf_net364));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net873 (.A(net873),
    .X(clknet_0_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net873 (.A(clknet_0_net873),
    .X(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net873 (.A(clknet_0_net873),
    .X(clknet_1_1__leaf_net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net899 (.A(net899),
    .X(clknet_0_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net171 (.A(net171),
    .X(clknet_0_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_0__leaf_net171));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net171 (.A(clknet_0_net171),
    .X(clknet_1_1__leaf_net171));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net14),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net938),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net939),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net881),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net941),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net22),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net943),
    .X(net944));
 sky130_fd_sc_hd__buf_2 rebuffer8 (.A(net943),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net887),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net946),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net389),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net948),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net662),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net950),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net887),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net152),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net954),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net389),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net662),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net895),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net253),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net751),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net704),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net772),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net727),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net698),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net707),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net732),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net464),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net564),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net239),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net777),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net859),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net430),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net251),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net865),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net778),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net703),
    .X(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A (.DIODE(net0));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1_N (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_Y (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A4 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_Y (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_Y (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1_N (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1_N (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_Y (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SET_B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCE (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_SET_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCD (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_RESET_B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A4 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_Y (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_SET_B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_SCE (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_D (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_SET_B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A4 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_RESET_B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_DE (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCE (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCE (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A4 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1_N (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_RESET_B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCD (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_Q (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_SET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A4 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A4 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A4 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A4 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B1_N (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q_N (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_RESET_B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A4 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_Q (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_Q_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCD (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCD (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A4 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_Q_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A4 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_Q (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_SCD (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A4 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B1_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_S1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_Y (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Y (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1_N (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Y (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_Y (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_S0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_Y (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCD (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A4 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SCD (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A4 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_RESET_B (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_B1_N (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_D (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_D (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_Q (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_X (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_X (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCD (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_Y (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net416_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SCE (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B1_N (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SCE (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q_N (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_Y (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q_N (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_Q_N (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_Q (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCE (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SCE (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCD (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_SCD (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_Y (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_Y (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_B1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_X (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_RESET_B (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_X (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_Y (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B1_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B1_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A4 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q_N (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A4 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1_N (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_Q (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCE (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_s833_Q (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_SET_B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_B1_N (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B1_N (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_SCE (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_Q (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B1_N (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_Q (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_SCE (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_Q_N (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCE (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SCE (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_Q (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A4 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q_N (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1_N (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1_N (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_Q (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A4 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A4 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_Q (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_Q_N (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_RESET_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCD (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_Y (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1_N (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_D (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_RESET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1_N (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1_N (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCE (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_RESET_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_D (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1_N (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_S1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_D (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_B1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_SET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1_N (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_RESET_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_Y (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S0 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_X (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_Q (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_Q_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_Q (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_SCD (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_Q (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_SCE (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_Q (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_Q (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCE (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_Q (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1_N (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A2 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_B1_N (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A4 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCE (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCD (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B1_N (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_D (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SCD (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_SCE (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B1_N (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1_N (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_DE (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SCD (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1_N (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_D (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B1_N (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B1_N (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_SCD (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCD (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SCE (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_SET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B1_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B1_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B1_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1_N (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1_N (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A4 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SET_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_SET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_SLEEP_B (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s833_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B1_N (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A4 (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net407_X (.DIODE(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SET_B (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_D (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net407_X (.DIODE(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_SCE (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A4 (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net860_X (.DIODE(clknet_1_0__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SCD (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A4 (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net860_X (.DIODE(clknet_1_1__leaf_net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net861_X (.DIODE(clknet_1_1__leaf_net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SET_B (.DIODE(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net873_X (.DIODE(clknet_1_0__leaf_net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SET_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_X (.DIODE(net961));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net900),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_1 clone2 (.A(net900),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net1),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net38),
    .X(net980));
 sky130_fd_sc_hd__a41o_1 clone22 (.A1(net72),
    .A2(net73),
    .A3(net67),
    .A4(net64),
    .B1(net71),
    .X(net981));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
