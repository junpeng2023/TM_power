module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net422;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net808;
 wire clknet_1_0__leaf_net808;
 wire clknet_1_1__leaf_net808;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net614;
 wire clknet_1_0__leaf_net614;
 wire clknet_1_1__leaf_net614;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net582;
 wire clknet_1_0__leaf_net582;
 wire clknet_1_1__leaf_net582;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net610;
 wire clknet_1_0__leaf_net610;
 wire clknet_1_1__leaf_net610;
 wire clknet_0_net624;
 wire clknet_1_0__leaf_net624;
 wire clknet_1_1__leaf_net624;
 wire clknet_0_net642;
 wire clknet_1_0__leaf_net642;
 wire clknet_1_1__leaf_net642;
 wire clknet_0_net643;
 wire clknet_1_0__leaf_net643;
 wire clknet_1_1__leaf_net643;
 wire clknet_0_net807;
 wire clknet_1_0__leaf_net807;
 wire clknet_1_1__leaf_net807;
 wire clknet_0_net806;
 wire clknet_1_0__leaf_net806;
 wire clknet_1_1__leaf_net806;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net512;
 wire clknet_1_0__leaf_net512;
 wire clknet_1_1__leaf_net512;
 wire clknet_0_net511;
 wire clknet_1_0__leaf_net511;
 wire clknet_1_1__leaf_net511;
 wire clknet_0_net790;
 wire clknet_1_0__leaf_net790;
 wire clknet_1_1__leaf_net790;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net789;
 wire clknet_1_0__leaf_net789;
 wire clknet_1_1__leaf_net789;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net741;
 wire clknet_1_0__leaf_net741;
 wire clknet_1_1__leaf_net741;
 wire clknet_0_net907;
 wire clknet_1_0__leaf_net907;
 wire clknet_1_1__leaf_net907;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net908;
 wire clknet_1_0__leaf_net908;
 wire clknet_1_1__leaf_net908;
 wire clknet_0_net277;
 wire clknet_1_0__leaf_net277;
 wire clknet_1_1__leaf_net277;
 wire clknet_0_net770;
 wire clknet_1_0__leaf_net770;
 wire clknet_1_1__leaf_net770;
 wire clknet_0_net508;
 wire clknet_1_0__leaf_net508;
 wire clknet_1_1__leaf_net508;
 wire clknet_0_net628;
 wire clknet_1_0__leaf_net628;
 wire clknet_1_1__leaf_net628;
 wire clknet_0_net930;
 wire clknet_1_0__leaf_net930;
 wire clknet_1_1__leaf_net930;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire clknet_0_net524;
 wire clknet_1_0__leaf_net524;
 wire clknet_1_1__leaf_net524;
 wire clknet_0_net263;
 wire clknet_1_0__leaf_net263;
 wire clknet_1_1__leaf_net263;
 wire clknet_0_net285;
 wire clknet_1_0__leaf_net285;
 wire clknet_1_1__leaf_net285;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net288;
 wire clknet_1_0__leaf_net288;
 wire clknet_1_1__leaf_net288;
 wire clknet_0_net284;
 wire clknet_1_0__leaf_net284;
 wire clknet_1_1__leaf_net284;
 wire clknet_0_net768;
 wire clknet_1_0__leaf_net768;
 wire clknet_1_1__leaf_net768;
 wire clknet_0_net275;
 wire clknet_1_0__leaf_net275;
 wire clknet_1_1__leaf_net275;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net63;
 wire clknet_1_0__leaf_net63;
 wire clknet_1_1__leaf_net63;
 wire clknet_0_net267;
 wire clknet_1_0__leaf_net267;
 wire clknet_1_1__leaf_net267;
 wire clknet_0_net928;
 wire clknet_1_0__leaf_net928;
 wire clknet_1_1__leaf_net928;
 wire clknet_0_net415;
 wire clknet_1_0__leaf_net415;
 wire clknet_1_1__leaf_net415;
 wire clknet_0_net400;
 wire clknet_1_0__leaf_net400;
 wire clknet_1_1__leaf_net400;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net252;
 wire clknet_1_0__leaf_net252;
 wire clknet_1_1__leaf_net252;
 wire clknet_0_net253;
 wire clknet_1_0__leaf_net253;
 wire clknet_1_1__leaf_net253;
 wire clknet_0_net264;
 wire clknet_1_0__leaf_net264;
 wire clknet_1_1__leaf_net264;
 wire clknet_0_net740;
 wire clknet_1_0__leaf_net740;
 wire clknet_1_1__leaf_net740;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net916;
 wire clknet_1_0__leaf_net916;
 wire clknet_1_1__leaf_net916;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net913;
 wire clknet_1_0__leaf_net913;
 wire clknet_1_1__leaf_net913;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net152;
 wire clknet_1_0__leaf_net152;
 wire clknet_1_1__leaf_net152;
 wire clknet_0_net281;
 wire clknet_1_0__leaf_net281;
 wire clknet_1_1__leaf_net281;
 wire clknet_0_net880;
 wire clknet_1_0__leaf_net880;
 wire clknet_1_1__leaf_net880;
 wire clknet_0_net173;
 wire clknet_1_0__leaf_net173;
 wire clknet_1_1__leaf_net173;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire clknet_0_net151;
 wire clknet_1_0__leaf_net151;
 wire clknet_1_1__leaf_net151;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;

 sky130_fd_sc_hd__or4bb_4 c100 (.A(net26),
    .B(net872),
    .C_N(net22),
    .D_N(net33),
    .X(net37));
 sky130_fd_sc_hd__and3_1 c101 (.A(net30),
    .B(net13),
    .C(net34),
    .X(net38));
 sky130_fd_sc_hd__and3_1 c102 (.A(net35),
    .B(net962),
    .C(net37),
    .X(net39));
 sky130_fd_sc_hd__and3_1 c103 (.A(net34),
    .B(net31),
    .C(net26),
    .X(net40));
 sky130_fd_sc_hd__and2_1 c104 (.A(net40),
    .B(net35),
    .X(net41));
 sky130_fd_sc_hd__and2_2 c105 (.A(net36),
    .B(net39),
    .X(net923));
 sky130_fd_sc_hd__or4bb_1 c106 (.A(net859),
    .B(net33),
    .C_N(net38),
    .D_N(net923),
    .X(net42));
 sky130_fd_sc_hd__and3_1 c107 (.A(net38),
    .B(net41),
    .C(net691),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 c108 (.A(net994),
    .X(net44));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net33),
    .A1(net44),
    .A2(net962),
    .A3(net43),
    .S0(net35),
    .S1(net31),
    .X(net45));
 sky130_fd_sc_hd__and2_0 c110 (.A(net843),
    .B(net826),
    .X(net46));
 sky130_fd_sc_hd__and2_0 c111 (.A(net28),
    .B(net826),
    .X(net47));
 sky130_fd_sc_hd__and2_0 c112 (.A(net25),
    .B(net28),
    .X(net48));
 sky130_fd_sc_hd__and2_1 c113 (.A(net852),
    .B(net2),
    .X(net49));
 sky130_fd_sc_hd__and2_0 c114 (.A(net826),
    .B(net31),
    .X(net50));
 sky130_fd_sc_hd__a2111o_1 c115 (.A1(net2),
    .A2(net944),
    .B1(net50),
    .C1(net37),
    .D1(net28),
    .X(net51));
 sky130_fd_sc_hd__and3_2 c116 (.A(net51),
    .B(net962),
    .C(net870),
    .X(net52));
 sky130_fd_sc_hd__and2_1 c117 (.A(net858),
    .B(net13),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c118 (.A(net46),
    .B(net53),
    .X(net54));
 sky130_fd_sc_hd__and2_1 c119 (.A(net46),
    .B(net52),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 c120 (.A(net761),
    .X(net915));
 sky130_fd_sc_hd__and3_1 c121 (.A(net50),
    .B(net944),
    .C(net53),
    .X(net56));
 sky130_fd_sc_hd__sdfbbn_1 c122 (.CLK_N(clknet_4_15_0_clk),
    .D(net56),
    .RESET_B(net55),
    .SCD(net49),
    .SCE(net53),
    .SET_B(net31),
    .Q(net884),
    .Q_N(net57));
 sky130_fd_sc_hd__and3_1 c123 (.A(net56),
    .B(net884),
    .C(net13),
    .X(net58));
 sky130_fd_sc_hd__buf_2 c124 (.A(net761),
    .X(net917));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net13),
    .A1(net47),
    .A2(net51),
    .A3(net25),
    .S0(net52),
    .S1(net57),
    .X(net59));
 sky130_fd_sc_hd__a2111o_1 c126 (.A1(net58),
    .A2(net49),
    .B1(net59),
    .C1(net2),
    .D1(net52),
    .X(net60));
 sky130_fd_sc_hd__mux4_1 c127 (.A0(net49),
    .A1(net884),
    .A2(net59),
    .A3(net13),
    .S0(net52),
    .S1(net25),
    .X(net61));
 sky130_fd_sc_hd__and3_1 c128 (.A(net39),
    .B(net917),
    .C(net52),
    .X(net62));
 sky130_fd_sc_hd__and3_1 c129 (.A(net962),
    .B(net53),
    .C(clknet_1_1__leaf_net769),
    .X(net63));
 sky130_fd_sc_hd__sdfrbp_1 c130 (.CLK(clknet_4_15_0_clk),
    .D(net62),
    .RESET_B(clknet_1_0__leaf_net63),
    .SCD(net13),
    .SCE(net49),
    .Q(net927),
    .Q_N(net64));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net48),
    .A1(clknet_1_1__leaf_net63),
    .A2(net62),
    .A3(net843),
    .S0(net57),
    .S1(net55),
    .X(net65));
 sky130_fd_sc_hd__and3_1 c132 (.A(net820),
    .B(net863),
    .C(net877),
    .X(net66));
 sky130_fd_sc_hd__and3_1 c133 (.A(net831),
    .B(net422),
    .C(net830),
    .X(net67));
 sky130_fd_sc_hd__and2_0 c134 (.A(net67),
    .B(net66),
    .X(net68));
 sky130_fd_sc_hd__or4bb_1 c135 (.A(net422),
    .B(net68),
    .C_N(net863),
    .D_N(net832),
    .X(net69));
 sky130_fd_sc_hd__and2_1 c136 (.A(net832),
    .B(net67),
    .X(net70));
 sky130_fd_sc_hd__and2_4 c137 (.A(net863),
    .B(net67),
    .X(net71));
 sky130_fd_sc_hd__and2_1 c138 (.A(net68),
    .B(net827),
    .X(net72));
 sky130_fd_sc_hd__or4bb_1 c139 (.A(net71),
    .B(net820),
    .C_N(net877),
    .D_N(net67),
    .X(net73));
 sky130_fd_sc_hd__and2_4 c140 (.A(net821),
    .B(net73),
    .X(net74));
 sky130_fd_sc_hd__a2111o_4 c141 (.A1(net72),
    .A2(net830),
    .B1(net831),
    .C1(net827),
    .D1(net71),
    .X(net906));
 sky130_fd_sc_hd__and2_1 c142 (.A(net830),
    .B(net832),
    .X(net75));
 sky130_fd_sc_hd__and3_1 c143 (.A(net829),
    .B(net75),
    .C(net823),
    .X(net76));
 sky130_fd_sc_hd__and2_2 c144 (.A(net879),
    .B(net68),
    .X(net77));
 sky130_fd_sc_hd__a2111o_1 c145 (.A1(net76),
    .A2(net841),
    .B1(net422),
    .C1(net67),
    .D1(net831),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c146 (.A(net73),
    .B(net822),
    .X(net79));
 sky130_fd_sc_hd__and2_2 c147 (.A(net877),
    .B(net823),
    .X(net80));
 sky130_fd_sc_hd__or4bb_1 c148 (.A(net75),
    .B(net827),
    .C_N(net80),
    .D_N(net77),
    .X(net81));
 sky130_fd_sc_hd__and2_4 c149 (.A(net78),
    .B(net79),
    .X(net82));
 sky130_fd_sc_hd__and3_2 c150 (.A(net82),
    .B(net77),
    .C(net78),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net77),
    .A1(net83),
    .A2(net70),
    .A3(net80),
    .S0(net832),
    .S1(net74),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net66),
    .A1(net79),
    .A2(net81),
    .A3(net72),
    .S0(net829),
    .S1(net78),
    .X(net85));
 sky130_fd_sc_hd__a2111o_1 c153 (.A1(net69),
    .A2(net83),
    .B1(net820),
    .C1(net79),
    .D1(net82),
    .X(net86));
 sky130_fd_sc_hd__and3_4 c154 (.A(net819),
    .B(net846),
    .C(net847),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c155 (.A(net841),
    .B(net989),
    .X(net88));
 sky130_fd_sc_hd__and2_1 c156 (.A(net843),
    .B(net827),
    .X(net89));
 sky130_fd_sc_hd__and2_0 c157 (.A(net853),
    .B(net836),
    .X(net90));
 sky130_fd_sc_hd__and3_4 c158 (.A(net958),
    .B(net89),
    .C(net854),
    .X(net91));
 sky130_fd_sc_hd__and3_1 c159 (.A(net91),
    .B(net819),
    .C(net958),
    .X(net92));
 sky130_fd_sc_hd__and3_1 c160 (.A(net89),
    .B(net833),
    .C(net989),
    .X(net93));
 sky130_fd_sc_hd__and2_1 c161 (.A(net856),
    .B(net836),
    .X(net94));
 sky130_fd_sc_hd__and2_1 c162 (.A(net93),
    .B(net1021),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net94),
    .A1(net834),
    .A2(net90),
    .A3(net846),
    .S0(net833),
    .S1(net958),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c164 (.A(net91),
    .B(net90),
    .C(net80),
    .X(net97));
 sky130_fd_sc_hd__or4bb_4 c165 (.A(net97),
    .B(net846),
    .C_N(net839),
    .D_N(net959),
    .X(net98));
 sky130_fd_sc_hd__and2_4 c166 (.A(net98),
    .B(net92),
    .X(net99));
 sky130_fd_sc_hd__and2_1 c167 (.A(net98),
    .B(net89),
    .X(net100));
 sky130_fd_sc_hd__and3_4 c168 (.A(net100),
    .B(net94),
    .C(net958),
    .X(net101));
 sky130_fd_sc_hd__or4bb_4 c169 (.A(net94),
    .B(net99),
    .C_N(net100),
    .D_N(net958),
    .X(net102));
 sky130_fd_sc_hd__and3_1 c170 (.A(net102),
    .B(net89),
    .C(net97),
    .X(net103));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net70),
    .A1(net102),
    .A2(net99),
    .A3(net89),
    .S0(net82),
    .S1(net101),
    .X(net104));
 sky130_fd_sc_hd__and3_1 c172 (.A(net79),
    .B(net96),
    .C(net94),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c173 (.A0(net96),
    .A1(net100),
    .A2(net98),
    .A3(net94),
    .S0(net848),
    .S1(net105),
    .X(net106));
 sky130_fd_sc_hd__or4bb_4 c174 (.A(net104),
    .B(net841),
    .C_N(net103),
    .D_N(net989),
    .X(net107));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net107),
    .A1(net104),
    .A2(net92),
    .A3(net83),
    .S0(net91),
    .S1(net101),
    .X(net108));
 sky130_fd_sc_hd__and2_2 c176 (.A(net838),
    .B(net829),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c177 (.A(net3),
    .B(net91),
    .X(net110));
 sky130_fd_sc_hd__or4bb_4 c178 (.A(net857),
    .B(net865),
    .C_N(net106),
    .D_N(net108),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c179 (.A(net108),
    .B(net871),
    .C(net840),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c180 (.A(net864),
    .B(net966),
    .C(net872),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c181 (.A(net834),
    .B(net80),
    .C(net990),
    .X(net114));
 sky130_fd_sc_hd__and2_1 c182 (.A(net847),
    .B(net872),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c183 (.A(net819),
    .B(net857),
    .C(net990),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c184 (.A(net872),
    .B(net105),
    .C(net80),
    .X(net117));
 sky130_fd_sc_hd__and3_4 c185 (.A(net81),
    .B(net91),
    .C(net113),
    .X(net118));
 sky130_fd_sc_hd__and3_4 c186 (.A(net112),
    .B(net862),
    .C(net959),
    .X(net889));
 sky130_fd_sc_hd__and3_1 c187 (.A(net865),
    .B(net889),
    .C(net117),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(net105),
    .A1(net967),
    .A2(net115),
    .A3(net119),
    .S0(net961),
    .S1(net83),
    .X(net120));
 sky130_fd_sc_hd__or4bb_4 c189 (.A(net966),
    .B(net101),
    .C_N(net871),
    .D_N(net118),
    .X(net896));
 sky130_fd_sc_hd__or4bb_4 c190 (.A(net83),
    .B(net889),
    .C_N(net115),
    .D_N(net1),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c191 (.A0(net117),
    .A1(net1),
    .A2(net95),
    .A3(net121),
    .S0(net115),
    .S1(net862),
    .X(net122));
 sky130_fd_sc_hd__and3_1 c192 (.A(net122),
    .B(net117),
    .C(net105),
    .X(net123));
 sky130_fd_sc_hd__and3_2 c193 (.A(net119),
    .B(net106),
    .C(net118),
    .X(net124));
 sky130_fd_sc_hd__mux4_2 c194 (.A0(net115),
    .A1(net123),
    .A2(net119),
    .A3(net121),
    .S0(net971),
    .S1(net122),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net835),
    .A1(net3),
    .A2(net125),
    .A3(net981),
    .S0(net114),
    .S1(net990),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 c196 (.A(net709),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net123),
    .A1(net127),
    .A2(net117),
    .A3(net1),
    .S0(net124),
    .S1(clknet_1_1__leaf_net740),
    .X(net128));
 sky130_fd_sc_hd__and3_1 c198 (.A(net110),
    .B(net111),
    .C(clknet_1_1__leaf_net740),
    .X(net129));
 sky130_fd_sc_hd__mux4_2 c199 (.A0(net20),
    .A1(net896),
    .A2(net10),
    .A3(net7),
    .S0(net101),
    .S1(net959),
    .X(net130));
 sky130_fd_sc_hd__and3_1 c200 (.A(net106),
    .B(net124),
    .C(net108),
    .X(net131));
 sky130_fd_sc_hd__and3_2 c201 (.A(net827),
    .B(net861),
    .C(net824),
    .X(net132));
 sky130_fd_sc_hd__and3_1 c202 (.A(net15),
    .B(net118),
    .C(net130),
    .X(net133));
 sky130_fd_sc_hd__and3_4 c203 (.A(net130),
    .B(net110),
    .C(net15),
    .X(net134));
 sky130_fd_sc_hd__and3_2 c204 (.A(net844),
    .B(net71),
    .C(net15),
    .X(net135));
 sky130_fd_sc_hd__and3_1 c205 (.A(net860),
    .B(net101),
    .C(net110),
    .X(net136));
 sky130_fd_sc_hd__or4bb_1 c206 (.A(net10),
    .B(net833),
    .C_N(net132),
    .D_N(net133),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 c207 (.A(net774),
    .X(net138));
 sky130_fd_sc_hd__and3_1 c208 (.A(net130),
    .B(net20),
    .C(net990),
    .X(net139));
 sky130_fd_sc_hd__or4bb_1 c209 (.A(net24),
    .B(net826),
    .C_N(net139),
    .D_N(net774),
    .X(net140));
 sky130_fd_sc_hd__buf_1 c210 (.A(net774),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net136),
    .A1(net141),
    .A2(net132),
    .A3(net17),
    .S0(net983),
    .S1(net962),
    .X(net142));
 sky130_fd_sc_hd__and3_1 c212 (.A(clknet_1_0__leaf_net129),
    .B(net111),
    .C(net136),
    .X(net143));
 sky130_fd_sc_hd__and3_1 c213 (.A(net871),
    .B(net136),
    .C(clknet_1_0__leaf_net143),
    .X(net144));
 sky130_fd_sc_hd__and3_1 c214 (.A(net17),
    .B(net130),
    .C(clknet_1_1__leaf_net740),
    .X(net145));
 sky130_fd_sc_hd__and3_1 c215 (.A(net131),
    .B(clknet_1_0__leaf_net143),
    .C(net136),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net133),
    .A1(net130),
    .A2(net134),
    .A3(clknet_1_0__leaf_net145),
    .S0(clknet_1_1__leaf_net129),
    .S1(net141),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net146),
    .A1(clknet_1_0__leaf_net144),
    .A2(clknet_1_1__leaf_net145),
    .A3(net1021),
    .S0(net141),
    .S1(net783),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(clknet_1_0__leaf_net145),
    .A1(net136),
    .A2(net20),
    .A3(net10),
    .S0(net141),
    .S1(net783),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net138),
    .A1(net134),
    .A2(net774),
    .A3(net782),
    .S0(net784),
    .S1(net786),
    .X(net150));
 sky130_fd_sc_hd__and3_4 c220 (.A(net34),
    .B(net7),
    .C(net961),
    .X(net901));
 sky130_fd_sc_hd__and3_1 c221 (.A(net968),
    .B(net37),
    .C(clknet_1_0__leaf_net144),
    .X(net151));
 sky130_fd_sc_hd__and2_0 c222 (.A(net44),
    .B(clknet_1_1__leaf_net143),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net994),
    .X(net153));
 sky130_fd_sc_hd__and3_1 c224 (.A(net17),
    .B(net101),
    .C(net98),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net41),
    .A1(net944),
    .A2(net923),
    .A3(net858),
    .S0(net34),
    .S1(net785),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c226 (.A(net136),
    .B(clknet_1_1__leaf_net152),
    .C(net691),
    .X(net156));
 sky130_fd_sc_hd__and3_1 c227 (.A(net154),
    .B(net34),
    .C(net71),
    .X(net157));
 sky130_fd_sc_hd__and3_1 c228 (.A(clknet_1_0__leaf_net156),
    .B(net37),
    .C(net154),
    .X(net158));
 sky130_fd_sc_hd__and3_1 c229 (.A(net153),
    .B(net135),
    .C(net17),
    .X(net159));
 sky130_fd_sc_hd__and3_1 c230 (.A(net159),
    .B(clknet_1_1__leaf_net156),
    .C(net154),
    .X(net160));
 sky130_fd_sc_hd__or4bb_4 c231 (.A(net833),
    .B(net41),
    .C_N(net872),
    .D_N(net783),
    .X(net161));
 sky130_fd_sc_hd__or4bb_1 c232 (.A(clknet_1_0__leaf_net156),
    .B(net828),
    .C_N(clknet_1_1__leaf_net143),
    .D_N(net154),
    .X(net162));
 sky130_fd_sc_hd__sdfrbp_1 c233 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net162),
    .RESET_B(net153),
    .SCD(net159),
    .SCE(net157),
    .Q(net164),
    .Q_N(net163));
 sky130_fd_sc_hd__sdfbbn_1 c234 (.CLK_N(clknet_4_15_0_clk),
    .D(net160),
    .RESET_B(net985),
    .SCD(net164),
    .SCE(net157),
    .SET_B(net691),
    .Q(net166),
    .Q_N(net165));
 sky130_fd_sc_hd__and3_2 c235 (.A(net861),
    .B(net164),
    .C(net157),
    .X(net167));
 sky130_fd_sc_hd__or4bb_1 c236 (.A(clknet_1_1__leaf_net158),
    .B(clknet_1_1__leaf_net162),
    .C_N(net159),
    .D_N(net167),
    .X(net168));
 sky130_fd_sc_hd__a2111o_1 c237 (.A1(net166),
    .A2(net135),
    .B1(net163),
    .C1(net734),
    .D1(net785),
    .X(net169));
 sky130_fd_sc_hd__sdfbbp_1 c238 (.CLK(clknet_4_13_0_clk),
    .D(net134),
    .RESET_B(net968),
    .SCD(net161),
    .SCE(clknet_1_0__leaf_net143),
    .SET_B(net167),
    .Q(net171),
    .Q_N(net170));
 sky130_fd_sc_hd__a2111o_1 c239 (.A1(net166),
    .A2(net167),
    .B1(net159),
    .C1(net972),
    .D1(net994),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net157),
    .A1(clknet_1_1__leaf_net152),
    .A2(net169),
    .A3(net163),
    .S0(clknet_1_1__leaf_net156),
    .S1(net167),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net872),
    .A1(net169),
    .A2(clknet_1_0__leaf_net158),
    .A3(net25),
    .S0(clknet_1_1__leaf_net152),
    .S1(net784),
    .X(net174));
 sky130_fd_sc_hd__and3_1 c242 (.A(net121),
    .B(net843),
    .C(clknet_1_1__leaf_net143),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c243 (.A(clknet_1_1__leaf_net143),
    .B(net944),
    .C(net901),
    .X(net176));
 sky130_fd_sc_hd__and3_1 c244 (.A(net47),
    .B(net962),
    .C(net897),
    .X(net177));
 sky130_fd_sc_hd__and3_2 c245 (.A(net47),
    .B(net54),
    .C(net901),
    .X(net178));
 sky130_fd_sc_hd__or4bb_1 c246 (.A(net53),
    .B(clknet_1_1__leaf_net144),
    .C_N(net167),
    .D_N(clknet_1_1__leaf_net175),
    .X(net913));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(clknet_1_1__leaf_net144),
    .A1(net25),
    .A2(net118),
    .A3(net52),
    .S0(clknet_1_0__leaf_net175),
    .S1(net917),
    .X(net179));
 sky130_fd_sc_hd__and3_1 c248 (.A(net58),
    .B(net962),
    .C(net843),
    .X(net180));
 sky130_fd_sc_hd__and3_1 c249 (.A(net176),
    .B(net927),
    .C(net167),
    .X(net916));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(clknet_1_0__leaf_net175),
    .A1(net52),
    .A2(net944),
    .A3(net55),
    .S0(net121),
    .S1(net167),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 c251 (.A(net758),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c252 (.A0(net52),
    .A1(net178),
    .A2(net167),
    .A3(net977),
    .S0(net161),
    .S1(net985),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net182),
    .A1(net901),
    .A2(clknet_1_1__leaf_net144),
    .A3(clknet_1_1__leaf_net179),
    .S0(net180),
    .S1(net787),
    .X(net184));
 sky130_fd_sc_hd__and3_1 c254 (.A(net180),
    .B(net781),
    .C(net787),
    .X(net185));
 sky130_fd_sc_hd__and3_1 c255 (.A(net185),
    .B(net167),
    .C(net759),
    .X(net186));
 sky130_fd_sc_hd__a2111o_1 c256 (.A1(net101),
    .A2(clknet_1_1__leaf_net179),
    .B1(net185),
    .C1(net177),
    .D1(net178),
    .X(net187));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net80),
    .A1(net182),
    .A2(net177),
    .A3(net31),
    .S0(net962),
    .S1(clknet_1_1__leaf_net179),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net866),
    .A1(net101),
    .A2(clknet_1_1__leaf_net179),
    .A3(net739),
    .S0(net781),
    .S1(net788),
    .X(net189));
 sky130_fd_sc_hd__mux4_2 c259 (.A0(net875),
    .A1(net31),
    .A2(net28),
    .A3(net178),
    .S0(net781),
    .S1(net788),
    .X(net190));
 sky130_fd_sc_hd__buf_1 c260 (.A(net758),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net191),
    .A1(net826),
    .A2(net190),
    .A3(clknet_1_0__leaf_net179),
    .S0(net739),
    .S1(net788),
    .X(net192));
 sky130_fd_sc_hd__buf_1 c262 (.A(clknet_1_1__leaf_net741),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net186),
    .A1(net190),
    .A2(net161),
    .A3(clknet_1_0__leaf_net179),
    .S0(net917),
    .S1(clknet_1_1__leaf_net741),
    .X(net194));
 sky130_fd_sc_hd__and2_1 c264 (.A(net75),
    .B(net76),
    .X(net195));
 sky130_fd_sc_hd__and2_1 c265 (.A(net86),
    .B(net74),
    .X(net196));
 sky130_fd_sc_hd__and2_2 c266 (.A(net74),
    .B(net76),
    .X(net197));
 sky130_fd_sc_hd__and2_2 c267 (.A(net826),
    .B(net82),
    .X(net198));
 sky130_fd_sc_hd__and2_2 c268 (.A(net86),
    .B(net197),
    .X(net199));
 sky130_fd_sc_hd__and2_4 c269 (.A(net824),
    .B(net198),
    .X(net200));
 sky130_fd_sc_hd__a2111o_1 c270 (.A1(net198),
    .A2(net197),
    .B1(net196),
    .C1(net85),
    .D1(net77),
    .X(net201));
 sky130_fd_sc_hd__and2_2 c271 (.A(net201),
    .B(net200),
    .X(net202));
 sky130_fd_sc_hd__and3_1 c272 (.A(net823),
    .B(net82),
    .C(net199),
    .X(net203));
 sky130_fd_sc_hd__and3_1 c273 (.A(net201),
    .B(net202),
    .C(net941),
    .X(net204));
 sky130_fd_sc_hd__or4bb_1 c274 (.A(net852),
    .B(net824),
    .C_N(net75),
    .D_N(net197),
    .X(net205));
 sky130_fd_sc_hd__and2_2 c275 (.A(net878),
    .B(net75),
    .X(net206));
 sky130_fd_sc_hd__and2_1 c276 (.A(net199),
    .B(net832),
    .X(net922));
 sky130_fd_sc_hd__and2_1 c277 (.A(net202),
    .B(net201),
    .X(net207));
 sky130_fd_sc_hd__a2111o_1 c278 (.A1(net207),
    .A2(net195),
    .B1(net945),
    .C1(net86),
    .D1(net82),
    .X(net208));
 sky130_fd_sc_hd__and2_4 c279 (.A(net205),
    .B(net207),
    .X(net914));
 sky130_fd_sc_hd__a2111o_2 c280 (.A1(net195),
    .A2(net208),
    .B1(net940),
    .C1(net945),
    .D1(net207),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c281 (.A(net209),
    .B(net76),
    .C(net207),
    .X(net210));
 sky130_fd_sc_hd__a2111o_1 c282 (.A1(net210),
    .A2(net198),
    .B1(net209),
    .C1(net206),
    .D1(net202),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net196),
    .A1(net211),
    .A2(net210),
    .A3(net206),
    .S0(net209),
    .S1(net198),
    .X(net212));
 sky130_fd_sc_hd__a2111o_1 c284 (.A1(net211),
    .A2(net210),
    .B1(net914),
    .C1(net941),
    .D1(net952),
    .X(net213));
 sky130_fd_sc_hd__or4bb_1 c285 (.A(net74),
    .B(net82),
    .C_N(net914),
    .D_N(net952),
    .X(net214));
 sky130_fd_sc_hd__and2_1 c286 (.A(net103),
    .B(net839),
    .X(net215));
 sky130_fd_sc_hd__and3_2 c287 (.A(net106),
    .B(net202),
    .C(net957),
    .X(net216));
 sky130_fd_sc_hd__and2_1 c288 (.A(net823),
    .B(net216),
    .X(net217));
 sky130_fd_sc_hd__and2_1 c289 (.A(net216),
    .B(net103),
    .X(net218));
 sky130_fd_sc_hd__and2_1 c290 (.A(net100),
    .B(net216),
    .X(net219));
 sky130_fd_sc_hd__and2_0 c291 (.A(net203),
    .B(net95),
    .X(net220));
 sky130_fd_sc_hd__a2111o_1 c292 (.A1(net218),
    .A2(net216),
    .B1(net88),
    .C1(net206),
    .D1(net957),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net214),
    .A1(net218),
    .A2(net197),
    .A3(net219),
    .S0(net100),
    .S1(net215),
    .X(net222));
 sky130_fd_sc_hd__and2_1 c294 (.A(net218),
    .B(net952),
    .X(net223));
 sky130_fd_sc_hd__and2_2 c295 (.A(net223),
    .B(net216),
    .X(net224));
 sky130_fd_sc_hd__and2_1 c296 (.A(net215),
    .B(net821),
    .X(net225));
 sky130_fd_sc_hd__and2_1 c297 (.A(net214),
    .B(net224),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 c298 (.A(net687),
    .X(net227));
 sky130_fd_sc_hd__or4bb_4 c299 (.A(net205),
    .B(net88),
    .C_N(net989),
    .D_N(net952),
    .X(net228));
 sky130_fd_sc_hd__and2_1 c300 (.A(net227),
    .B(net223),
    .X(net229));
 sky130_fd_sc_hd__and3_1 c301 (.A(net229),
    .B(net220),
    .C(net216),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c302 (.A(net222),
    .B(net217),
    .X(net231));
 sky130_fd_sc_hd__a2111o_1 c303 (.A1(net836),
    .A2(net230),
    .B1(net937),
    .C1(net989),
    .D1(net945),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net230),
    .A1(net839),
    .A2(net227),
    .A3(net214),
    .S0(net224),
    .S1(net226),
    .X(net233));
 sky130_fd_sc_hd__and3_1 c305 (.A(net103),
    .B(net229),
    .C(net952),
    .X(net234));
 sky130_fd_sc_hd__mux4_2 c306 (.A0(net229),
    .A1(net203),
    .A2(net108),
    .A3(net228),
    .S0(net223),
    .S1(net687),
    .X(net235));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net220),
    .A1(net227),
    .A2(net224),
    .A3(net197),
    .S0(net228),
    .S1(net687),
    .X(net236));
 sky130_fd_sc_hd__and2_1 c308 (.A(net228),
    .B(net120),
    .X(net237));
 sky130_fd_sc_hd__and2_2 c309 (.A(net205),
    .B(net237),
    .X(net238));
 sky130_fd_sc_hd__and3_1 c310 (.A(net114),
    .B(net228),
    .C(net71),
    .X(net239));
 sky130_fd_sc_hd__and2_1 c311 (.A(net223),
    .B(net108),
    .X(net240));
 sky130_fd_sc_hd__buf_1 c312 (.A(net767),
    .X(net241));
 sky130_fd_sc_hd__and2_0 c313 (.A(net95),
    .B(net961),
    .X(net242));
 sky130_fd_sc_hd__a2111o_4 c314 (.A1(net239),
    .A2(net219),
    .B1(net197),
    .C1(net223),
    .D1(net687),
    .X(net243));
 sky130_fd_sc_hd__and3_1 c315 (.A(net197),
    .B(net242),
    .C(net687),
    .X(net244));
 sky130_fd_sc_hd__buf_1 c316 (.A(net767),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c317 (.A(net869),
    .B(net108),
    .C(net85),
    .X(net246));
 sky130_fd_sc_hd__and3_1 c318 (.A(net120),
    .B(net240),
    .C(net245),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c319 (.A(net822),
    .B(net244),
    .C(net228),
    .X(net248));
 sky130_fd_sc_hd__mux4_2 c320 (.A0(net237),
    .A1(net246),
    .A2(net245),
    .A3(net200),
    .S0(net239),
    .S1(net240),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(net248),
    .A1(net914),
    .A2(net249),
    .A3(net237),
    .S0(net95),
    .S1(net199),
    .X(net250));
 sky130_fd_sc_hd__buf_1 c322 (.A(net767),
    .X(net251));
 sky130_fd_sc_hd__or4bb_1 c323 (.A(net219),
    .B(net111),
    .C_N(net985),
    .D_N(clknet_1_0__leaf_net789),
    .X(net252));
 sky130_fd_sc_hd__and3_1 c324 (.A(net242),
    .B(net239),
    .C(clknet_1_1__leaf_net252),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net245),
    .A1(net251),
    .A2(net197),
    .A3(net836),
    .S0(net243),
    .S1(net249),
    .X(net254));
 sky130_fd_sc_hd__a2111o_1 c326 (.A1(net246),
    .A2(net85),
    .B1(net241),
    .C1(net237),
    .D1(clknet_1_0__leaf_net790),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net240),
    .A1(net822),
    .A2(net251),
    .A3(net237),
    .S0(net243),
    .S1(clknet_1_1__leaf_net255),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(clknet_1_0__leaf_net255),
    .A1(net963),
    .A2(net121),
    .A3(net249),
    .S0(clknet_1_0__leaf_net789),
    .S1(clknet_1_0__leaf_net790),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net219),
    .A1(clknet_1_0__leaf_net255),
    .A2(net940),
    .A3(net216),
    .S0(net237),
    .S1(net767),
    .X(net258));
 sky130_fd_sc_hd__buf_1 c330 (.A(net752),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c331 (.A(net914),
    .B(net118),
    .C(net786),
    .X(net260));
 sky130_fd_sc_hd__or4bb_1 c332 (.A(net243),
    .B(net236),
    .C_N(net987),
    .D_N(clknet_1_0__leaf_net789),
    .X(net261));
 sky130_fd_sc_hd__and3_1 c333 (.A(net251),
    .B(net74),
    .C(net200),
    .X(net262));
 sky130_fd_sc_hd__and3_1 c334 (.A(net71),
    .B(net786),
    .C(clknet_1_1__leaf_net789),
    .X(net263));
 sky130_fd_sc_hd__and3_1 c335 (.A(clknet_1_0__leaf_net253),
    .B(net259),
    .C(net873),
    .X(net264));
 sky130_fd_sc_hd__sdfrtn_1 c336 (.CLK_N(clknet_4_12_0_clk),
    .D(net247),
    .RESET_B(net236),
    .SCD(clknet_1_0__leaf_net263),
    .SCE(clknet_1_0__leaf_net789),
    .Q(net265));
 sky130_fd_sc_hd__and3_1 c337 (.A(clknet_1_0__leaf_net252),
    .B(net940),
    .C(net873),
    .X(net266));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net858),
    .A1(net889),
    .A2(net828),
    .A3(clknet_1_0__leaf_net263),
    .S0(net265),
    .S1(net784),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net241),
    .A1(clknet_1_0__leaf_net267),
    .A2(net945),
    .A3(net231),
    .S0(net957),
    .S1(clknet_1_1__leaf_net789),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(net265),
    .A1(net259),
    .A2(net249),
    .A3(net135),
    .S0(clknet_1_1__leaf_net263),
    .S1(net961),
    .X(net269));
 sky130_fd_sc_hd__and3_1 c341 (.A(net260),
    .B(net132),
    .C(net786),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net259),
    .A1(net127),
    .A2(clknet_1_0__leaf_net263),
    .A3(net992),
    .S0(clknet_1_1__leaf_net253),
    .S1(net782),
    .X(net271));
 sky130_fd_sc_hd__and3_1 c343 (.A(net266),
    .B(net265),
    .C(net991),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net889),
    .A1(clknet_1_0__leaf_net264),
    .A2(clknet_1_0__leaf_net263),
    .A3(net270),
    .S0(net259),
    .S1(net767),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 c345 (.A(net752),
    .X(net274));
 sky130_fd_sc_hd__and3_1 c346 (.A(clknet_1_0__leaf_net267),
    .B(net127),
    .C(clknet_1_1__leaf_net768),
    .X(net275));
 sky130_fd_sc_hd__a2111o_1 c347 (.A1(clknet_1_0__leaf_net275),
    .A2(net265),
    .B1(net87),
    .C1(clknet_1_1__leaf_net768),
    .D1(clknet_1_1__leaf_net789),
    .X(net924));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net274),
    .A1(net970),
    .A2(clknet_1_0__leaf_net264),
    .A3(clknet_1_1__leaf_net275),
    .S0(net1016),
    .S1(net236),
    .X(net276));
 sky130_fd_sc_hd__or4bb_4 c349 (.A(net262),
    .B(clknet_1_0__leaf_net275),
    .C_N(clknet_1_0__leaf_net924),
    .D_N(net786),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net272),
    .A1(clknet_1_0__leaf_net275),
    .A2(net241),
    .A3(clknet_1_0__leaf_net277),
    .S0(net991),
    .S1(net767),
    .X(net278));
 sky130_fd_sc_hd__mux4_2 c351 (.A0(clknet_1_0__leaf_net275),
    .A1(clknet_1_1__leaf_net277),
    .A2(net265),
    .A3(net737),
    .S0(net767),
    .S1(clknet_1_0__leaf_net769),
    .X(net279));
 sky130_fd_sc_hd__and3_1 c352 (.A(net171),
    .B(net826),
    .C(clknet_1_0__leaf_net769),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(clknet_1_0__leaf_net152),
    .A1(net171),
    .A2(net118),
    .A3(net111),
    .S0(net31),
    .S1(net691),
    .X(net281));
 sky130_fd_sc_hd__and2_1 c354 (.A(net858),
    .B(net785),
    .X(net282));
 sky130_fd_sc_hd__or4bb_1 c355 (.A(net172),
    .B(clknet_1_1__leaf_net263),
    .C_N(clknet_1_1__leaf_net281),
    .D_N(net691),
    .X(net283));
 sky130_fd_sc_hd__and2_0 c356 (.A(net280),
    .B(clknet_1_1__leaf_net263),
    .X(net284));
 sky130_fd_sc_hd__and2_0 c357 (.A(net200),
    .B(clknet_1_1__leaf_net281),
    .X(net880));
 sky130_fd_sc_hd__and3_1 c358 (.A(clknet_1_1__leaf_net263),
    .B(clknet_1_0__leaf_net152),
    .C(clknet_1_0__leaf_net769),
    .X(net285));
 sky130_fd_sc_hd__sdfrtp_2 c359 (.CLK(clknet_4_14_0_clk),
    .D(net169),
    .RESET_B(net135),
    .SCD(clknet_1_1__leaf_net264),
    .SCE(clknet_1_1__leaf_net151),
    .Q(net286));
 sky130_fd_sc_hd__and3_1 c360 (.A(net169),
    .B(net940),
    .C(net774),
    .X(net287));
 sky130_fd_sc_hd__a2111o_1 c361 (.A1(clknet_1_1__leaf_net285),
    .A2(net961),
    .B1(net901),
    .C1(net170),
    .D1(net748),
    .X(net288));
 sky130_fd_sc_hd__and3_1 c362 (.A(clknet_1_0__leaf_net281),
    .B(clknet_1_0__leaf_net285),
    .C(clknet_1_1__leaf_net267),
    .X(net289));
 sky130_fd_sc_hd__buf_1 c363 (.A(clknet_1_1__leaf_net742),
    .X(net290));
 sky130_fd_sc_hd__sdfbbn_1 c364 (.CLK_N(clknet_4_12_0_clk),
    .D(net32),
    .RESET_B(clknet_1_1__leaf_net289),
    .SCD(net282),
    .SCE(net25),
    .SET_B(clknet_1_0__leaf_net281),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__or4bb_1 c365 (.A(net236),
    .B(net282),
    .C_N(net286),
    .D_N(clknet_1_1__leaf_net284),
    .X(net293));
 sky130_fd_sc_hd__buf_1 c366 (.A(clknet_1_1__leaf_net742),
    .X(net294));
 sky130_fd_sc_hd__a2111o_1 c367 (.A1(net1015),
    .A2(net291),
    .B1(clknet_1_0__leaf_net289),
    .C1(net747),
    .D1(clknet_1_0__leaf_net790),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net290),
    .A1(net292),
    .A2(clknet_1_0__leaf_net152),
    .A3(net910),
    .S0(clknet_1_1__leaf_net880),
    .S1(net774),
    .X(net296));
 sky130_fd_sc_hd__sdfbbn_1 c369 (.CLK_N(clknet_4_14_0_clk),
    .D(net1005),
    .RESET_B(net134),
    .SCD(net751),
    .SCE(net774),
    .SET_B(clknet_1_0__leaf_net931),
    .Q(net298),
    .Q_N(net297));
 sky130_fd_sc_hd__a2111o_1 c370 (.A1(net298),
    .A2(net292),
    .B1(clknet_1_1__leaf_net880),
    .C1(net286),
    .D1(net748),
    .X(net299));
 sky130_fd_sc_hd__a2111o_1 c371 (.A1(net292),
    .A2(net298),
    .B1(net691),
    .C1(net751),
    .D1(clknet_1_1__leaf_net790),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net287),
    .A1(net298),
    .A2(clknet_1_0__leaf_net300),
    .A3(net291),
    .S0(net946),
    .S1(net747),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(clknet_1_1__leaf_net300),
    .A1(net301),
    .A2(net200),
    .A3(net297),
    .S0(net972),
    .S1(clknet_1_0__leaf_net931),
    .X(net302));
 sky130_fd_sc_hd__or4bb_2 c374 (.A(net31),
    .B(net988),
    .C_N(net28),
    .D_N(net940),
    .X(net885));
 sky130_fd_sc_hd__or4bb_1 c375 (.A(net858),
    .B(net901),
    .C_N(net776),
    .D_N(net787),
    .X(net909));
 sky130_fd_sc_hd__and3_1 c376 (.A(net985),
    .B(net885),
    .C(clknet_1_1__leaf_net790),
    .X(net303));
 sky130_fd_sc_hd__sdfrtp_1 c377 (.CLK(clknet_4_14_0_clk),
    .D(net25),
    .RESET_B(net923),
    .SCD(net885),
    .SCE(net286),
    .Q(net304));
 sky130_fd_sc_hd__or4bb_2 c378 (.A(net286),
    .B(net884),
    .C_N(net987),
    .D_N(net748),
    .X(net918));
 sky130_fd_sc_hd__or4bb_2 c379 (.A(net178),
    .B(net917),
    .C_N(net64),
    .D_N(net177),
    .X(net903));
 sky130_fd_sc_hd__or4bb_1 c380 (.A(net161),
    .B(net855),
    .C_N(net944),
    .D_N(clknet_1_0__leaf_net741),
    .X(net305));
 sky130_fd_sc_hd__and3_1 c381 (.A(clknet_1_1__leaf_net193),
    .B(net918),
    .C(net748),
    .X(net898));
 sky130_fd_sc_hd__or4bb_1 c382 (.A(net304),
    .B(clknet_1_0__leaf_net916),
    .C_N(net914),
    .D_N(net178),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net55),
    .A1(net903),
    .A2(clknet_1_0__leaf_net193),
    .A3(net304),
    .S0(clknet_1_0__leaf_net179),
    .S1(clknet_1_1__leaf_net931),
    .X(net307));
 sky130_fd_sc_hd__a2111o_1 c384 (.A1(net191),
    .A2(net286),
    .B1(clknet_1_0__leaf_net179),
    .C1(net304),
    .D1(net761),
    .X(net308));
 sky130_fd_sc_hd__or4bb_1 c385 (.A(clknet_1_0__leaf_net179),
    .B(clknet_1_0__leaf_net898),
    .C_N(net191),
    .D_N(net914),
    .X(net309));
 sky130_fd_sc_hd__or4bb_1 c386 (.A(net177),
    .B(clknet_1_0__leaf_net898),
    .C_N(net918),
    .D_N(net921),
    .X(net920));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net178),
    .A1(net917),
    .A2(net37),
    .A3(clknet_1_0__leaf_net916),
    .S0(net886),
    .S1(clknet_1_1__leaf_net931),
    .X(net310));
 sky130_fd_sc_hd__sdfrtp_2 c388 (.CLK(clknet_4_14_0_clk),
    .D(net918),
    .RESET_B(net923),
    .SCD(net761),
    .SCE(clknet_1_1__leaf_net931),
    .Q(net311));
 sky130_fd_sc_hd__or4bb_1 c389 (.A(net118),
    .B(clknet_1_0__leaf_net913),
    .C_N(net311),
    .D_N(net787),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net303),
    .A1(net903),
    .A2(net311),
    .A3(net191),
    .S0(clknet_1_0__leaf_net916),
    .S1(net739),
    .X(net313));
 sky130_fd_sc_hd__or4bb_1 c391 (.A(net311),
    .B(net858),
    .C_N(net57),
    .D_N(net736),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net282),
    .A1(net161),
    .A2(net901),
    .A3(net311),
    .S0(net28),
    .S1(clknet_1_1__leaf_net790),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net54),
    .A1(clknet_1_1__leaf_net880),
    .A2(net311),
    .A3(net64),
    .S0(net918),
    .S1(net776),
    .X(net316));
 sky130_fd_sc_hd__a2111o_1 c394 (.A1(net191),
    .A2(net903),
    .B1(net945),
    .C1(net977),
    .D1(net776),
    .X(net317));
 sky130_fd_sc_hd__or4bb_1 c395 (.A(net314),
    .B(net311),
    .C_N(net739),
    .D_N(clknet_1_1__leaf_net769),
    .X(net929));
 sky130_fd_sc_hd__and2_1 c396 (.A(net67),
    .B(net84),
    .X(net318));
 sky130_fd_sc_hd__and2_1 c397 (.A(net825),
    .B(net204),
    .X(net319));
 sky130_fd_sc_hd__and2_2 c398 (.A(net85),
    .B(net942),
    .X(net320));
 sky130_fd_sc_hd__mux4_2 c399 (.A0(net74),
    .A1(net84),
    .A2(net825),
    .A3(net320),
    .S0(net942),
    .S1(net319),
    .X(net321));
 sky130_fd_sc_hd__and2_0 c400 (.A(net198),
    .B(net942),
    .X(net322));
 sky130_fd_sc_hd__and2_1 c401 (.A(net322),
    .B(net209),
    .X(net323));
 sky130_fd_sc_hd__and2_1 c402 (.A(net200),
    .B(net323),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c403 (.A0(net204),
    .A1(net324),
    .A2(net320),
    .A3(net318),
    .S0(net319),
    .S1(net323),
    .X(net325));
 sky130_fd_sc_hd__and2_2 c404 (.A(net321),
    .B(net952),
    .X(net326));
 sky130_fd_sc_hd__and2_1 c405 (.A(net323),
    .B(net326),
    .X(net327));
 sky130_fd_sc_hd__and2_1 c406 (.A(net77),
    .B(net682),
    .X(net328));
 sky130_fd_sc_hd__and2_1 c407 (.A(net328),
    .B(net320),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c408 (.A(net329),
    .B(net942),
    .C(net682),
    .X(net330));
 sky130_fd_sc_hd__buf_1 c409 (.A(net709),
    .X(net331));
 sky130_fd_sc_hd__and2_1 c410 (.A(net321),
    .B(net328),
    .X(net332));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(net321),
    .A1(net327),
    .A2(net319),
    .A3(net204),
    .S0(net942),
    .S1(net71),
    .X(net333));
 sky130_fd_sc_hd__and2_1 c412 (.A(net319),
    .B(net326),
    .X(net334));
 sky130_fd_sc_hd__buf_1 c413 (.A(net709),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net327),
    .A1(net321),
    .A2(net329),
    .A3(net332),
    .S0(net323),
    .S1(net198),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net334),
    .A1(net319),
    .A2(net330),
    .A3(net335),
    .S0(net320),
    .S1(net328),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net318),
    .A1(net331),
    .A2(net330),
    .A3(net321),
    .S0(net320),
    .S1(net794),
    .X(net338));
 sky130_fd_sc_hd__and3_1 c417 (.A(net338),
    .B(net335),
    .C(net320),
    .X(net339));
 sky130_fd_sc_hd__and2_1 c418 (.A(net850),
    .B(net940),
    .X(net340));
 sky130_fd_sc_hd__and2_2 c419 (.A(net202),
    .B(net88),
    .X(net902));
 sky130_fd_sc_hd__sdfbbp_1 c420 (.CLK(clknet_4_6_0_clk),
    .D(net334),
    .RESET_B(net945),
    .SCD(net226),
    .SCE(net957),
    .SET_B(net687),
    .Q(net887),
    .Q_N(net341));
 sky130_fd_sc_hd__and2_1 c421 (.A(net88),
    .B(net206),
    .X(net342));
 sky130_fd_sc_hd__and2_0 c422 (.A(net837),
    .B(net964),
    .X(net343));
 sky130_fd_sc_hd__buf_2 c423 (.A(net687),
    .X(net344));
 sky130_fd_sc_hd__and2_4 c424 (.A(net340),
    .B(net344),
    .X(net890));
 sky130_fd_sc_hd__a2111o_1 c425 (.A1(net331),
    .A2(net890),
    .B1(net839),
    .C1(net964),
    .D1(net955),
    .X(net345));
 sky130_fd_sc_hd__a2111o_1 c426 (.A1(net848),
    .A2(net821),
    .B1(net234),
    .C1(net217),
    .D1(net953),
    .X(net346));
 sky130_fd_sc_hd__and2_1 c427 (.A(net330),
    .B(net963),
    .X(net347));
 sky130_fd_sc_hd__or4bb_1 c428 (.A(net328),
    .B(net347),
    .C_N(net345),
    .D_N(net953),
    .X(net348));
 sky130_fd_sc_hd__and3_1 c429 (.A(net206),
    .B(net348),
    .C(net202),
    .X(net349));
 sky130_fd_sc_hd__mux4_2 c430 (.A0(net839),
    .A1(net206),
    .A2(net326),
    .A3(net963),
    .S0(net349),
    .S1(net684),
    .X(net350));
 sky130_fd_sc_hd__or4bb_4 c431 (.A(net217),
    .B(net955),
    .C_N(net348),
    .D_N(net224),
    .X(net351));
 sky130_fd_sc_hd__a2111o_1 c432 (.A1(net345),
    .A2(net351),
    .B1(net88),
    .C1(net953),
    .D1(net794),
    .X(net352));
 sky130_fd_sc_hd__a2111o_1 c433 (.A1(net329),
    .A2(net216),
    .B1(net942),
    .C1(net351),
    .D1(net953),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net335),
    .A1(net349),
    .A2(net340),
    .A3(net965),
    .S0(net342),
    .S1(net718),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net348),
    .A1(net354),
    .A2(net344),
    .A3(net226),
    .S0(net351),
    .S1(net791),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net343),
    .A1(net844),
    .A2(net350),
    .A3(net953),
    .S0(net683),
    .S1(net762),
    .X(net356));
 sky130_fd_sc_hd__or4bb_2 c437 (.A(net206),
    .B(net955),
    .C_N(net684),
    .D_N(net762),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net963),
    .A1(net235),
    .A2(net216),
    .A3(net351),
    .S0(net762),
    .S1(net1006),
    .X(net358));
 sky130_fd_sc_hd__a2111o_1 c439 (.A1(net354),
    .A2(net357),
    .B1(net206),
    .C1(net953),
    .D1(net763),
    .X(net359));
 sky130_fd_sc_hd__and2_0 c440 (.A(net961),
    .B(net199),
    .X(net360));
 sky130_fd_sc_hd__and2_0 c441 (.A(net957),
    .B(net794),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net244),
    .A1(net957),
    .A2(net344),
    .A3(net954),
    .S0(net687),
    .S1(net718),
    .X(net362));
 sky130_fd_sc_hd__and2_0 c443 (.A(net361),
    .B(net870),
    .X(net363));
 sky130_fd_sc_hd__sdfbbn_1 c444 (.CLK_N(clknet_4_6_0_clk),
    .D(net326),
    .RESET_B(net249),
    .SCD(net361),
    .SCE(net957),
    .SET_B(net953),
    .Q(net365),
    .Q_N(net364));
 sky130_fd_sc_hd__and2_1 c445 (.A(net868),
    .B(net342),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 c446 (.A(net709),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net360),
    .A1(net957),
    .A2(net367),
    .A3(net344),
    .S0(net200),
    .S1(net687),
    .X(net368));
 sky130_fd_sc_hd__and3_1 c448 (.A(net362),
    .B(net363),
    .C(net954),
    .X(net369));
 sky130_fd_sc_hd__a2111o_1 c449 (.A1(net1),
    .A2(net244),
    .B1(net364),
    .C1(net719),
    .D1(net793),
    .X(net370));
 sky130_fd_sc_hd__and3_1 c450 (.A(net113),
    .B(net365),
    .C(net326),
    .X(net371));
 sky130_fd_sc_hd__and2_2 c451 (.A(net216),
    .B(net360),
    .X(net372));
 sky130_fd_sc_hd__sdfbbn_1 c452 (.CLK_N(clknet_4_6_0_clk),
    .D(net368),
    .RESET_B(net999),
    .SCD(net74),
    .SCE(net957),
    .SET_B(net936),
    .Q(net374),
    .Q_N(net373));
 sky130_fd_sc_hd__a2111o_1 c453 (.A1(net344),
    .A2(net936),
    .B1(net326),
    .C1(net940),
    .D1(net754),
    .X(net375));
 sky130_fd_sc_hd__a2111o_1 c454 (.A1(net244),
    .A2(net121),
    .B1(net372),
    .C1(net326),
    .D1(net365),
    .X(net376));
 sky130_fd_sc_hd__sdfbbp_1 c455 (.CLK(clknet_4_6_0_clk),
    .D(net363),
    .RESET_B(net374),
    .SCD(net936),
    .SCE(net376),
    .SET_B(net762),
    .Q(net932),
    .Q_N(net377));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net365),
    .A1(net936),
    .A2(net326),
    .A3(net373),
    .S0(net868),
    .S1(net793),
    .X(net378));
 sky130_fd_sc_hd__sdfbbn_2 c457 (.CLK_N(clknet_4_9_0_clk),
    .D(net225),
    .RESET_B(net200),
    .SCD(net936),
    .SCE(net754),
    .SET_B(net1000),
    .Q(net380),
    .Q_N(net379));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net376),
    .A1(net373),
    .A2(net85),
    .A3(net380),
    .S0(net364),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net376),
    .A1(net344),
    .A2(net244),
    .A3(net957),
    .S0(net735),
    .S1(net754),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net351),
    .A1(net380),
    .A2(net936),
    .A3(net364),
    .S0(net687),
    .S1(net735),
    .X(net383));
 sky130_fd_sc_hd__sdfbbn_1 c461 (.CLK_N(clknet_4_6_0_clk),
    .D(net369),
    .RESET_B(net249),
    .SCD(net371),
    .SCE(net735),
    .SET_B(net795),
    .Q(net385),
    .Q_N(net384));
 sky130_fd_sc_hd__and2_1 c462 (.A(net367),
    .B(net763),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net270),
    .A1(net855),
    .A2(net231),
    .A3(net961),
    .S0(net954),
    .S1(net952),
    .X(net387));
 sky130_fd_sc_hd__and2_0 c464 (.A(net369),
    .B(net386),
    .X(net388));
 sky130_fd_sc_hd__buf_1 c465 (.A(clknet_1_1__leaf_net770),
    .X(net389));
 sky130_fd_sc_hd__and2_2 c466 (.A(net762),
    .B(net795),
    .X(net390));
 sky130_fd_sc_hd__and2_0 c467 (.A(net386),
    .B(net763),
    .X(net391));
 sky130_fd_sc_hd__and2_1 c468 (.A(net828),
    .B(net386),
    .X(net392));
 sky130_fd_sc_hd__and2_1 c469 (.A(net873),
    .B(net392),
    .X(net393));
 sky130_fd_sc_hd__sdfsbp_2 c470 (.CLK(clknet_4_9_0_clk),
    .D(net392),
    .SCD(net386),
    .SCE(net937),
    .SET_B(net995),
    .Q(net395),
    .Q_N(net394));
 sky130_fd_sc_hd__and2_0 c471 (.A(net370),
    .B(clknet_1_0__leaf_net742),
    .X(net396));
 sky130_fd_sc_hd__and2_0 c472 (.A(net395),
    .B(clknet_1_0__leaf_net768),
    .X(net397));
 sky130_fd_sc_hd__and3_1 c473 (.A(net395),
    .B(net852),
    .C(net738),
    .X(net398));
 sky130_fd_sc_hd__and2_1 c474 (.A(net392),
    .B(net796),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(net390),
    .A1(net393),
    .A2(net944),
    .A3(net391),
    .S0(clknet_1_0__leaf_net267),
    .S1(net796),
    .X(net400));
 sky130_fd_sc_hd__a2111o_1 c476 (.A1(net396),
    .A2(net399),
    .B1(net975),
    .C1(net372),
    .D1(net995),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net397),
    .A1(net399),
    .A2(net249),
    .A3(net852),
    .S0(net946),
    .S1(net961),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net391),
    .A1(net399),
    .A2(net844),
    .A3(net386),
    .S0(clknet_1_0__leaf_net400),
    .S1(net755),
    .X(net925));
 sky130_fd_sc_hd__a2111o_1 c479 (.A1(net389),
    .A2(net393),
    .B1(clknet_1_0__leaf_net925),
    .C1(net394),
    .D1(clknet_1_0__leaf_net742),
    .X(net930));
 sky130_fd_sc_hd__a2111o_1 c480 (.A1(net249),
    .A2(net393),
    .B1(net116),
    .C1(net1013),
    .D1(net797),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net393),
    .A1(clknet_1_1__leaf_net930),
    .A2(net249),
    .A3(clknet_1_0__leaf_net400),
    .S0(net394),
    .S1(net797),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net930),
    .A1(net380),
    .A2(net243),
    .A3(net399),
    .S0(net738),
    .S1(net797),
    .X(net405));
 sky130_fd_sc_hd__a2111o_1 c483 (.A1(net395),
    .A2(net367),
    .B1(net737),
    .C1(clknet_1_0__leaf_net768),
    .D1(net797),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(clknet_1_1__leaf_net288),
    .A1(net902),
    .A2(net200),
    .A3(net297),
    .S0(net398),
    .S1(clknet_1_0__leaf_net931),
    .X(net407));
 sky130_fd_sc_hd__a2111o_1 c485 (.A1(net401),
    .A2(net901),
    .B1(net890),
    .C1(clknet_1_0__leaf_net768),
    .D1(net798),
    .X(net408));
 sky130_fd_sc_hd__a2111o_1 c486 (.A1(net398),
    .A2(net225),
    .B1(net870),
    .C1(clknet_1_0__leaf_net925),
    .D1(net28),
    .X(net409));
 sky130_fd_sc_hd__and3_1 c487 (.A(net111),
    .B(clknet_1_1__leaf_net924),
    .C(clknet_1_0__leaf_net925),
    .X(net908));
 sky130_fd_sc_hd__a2111o_1 c488 (.A1(net225),
    .A2(net408),
    .B1(net828),
    .C1(clknet_1_1__leaf_net264),
    .D1(net798),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_4 c489 (.A(net752),
    .X(net411));
 sky130_fd_sc_hd__a2111o_1 c490 (.A1(net372),
    .A2(clknet_1_0__leaf_net924),
    .B1(net875),
    .C1(net783),
    .D1(net798),
    .X(net904));
 sky130_fd_sc_hd__a2111o_1 c491 (.A1(net28),
    .A2(clknet_1_0__leaf_net173),
    .B1(net411),
    .C1(clknet_1_0__leaf_net904),
    .D1(net946),
    .X(net412));
 sky130_fd_sc_hd__buf_1 c492 (.A(net752),
    .X(net413));
 sky130_fd_sc_hd__a2111o_1 c493 (.A1(net344),
    .A2(clknet_1_1__leaf_net880),
    .B1(net165),
    .C1(net875),
    .D1(net798),
    .X(net414));
 sky130_fd_sc_hd__a2111o_1 c494 (.A1(clknet_1_1__leaf_net267),
    .A2(net969),
    .B1(net691),
    .C1(net695),
    .D1(net798),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net388),
    .A1(net170),
    .A2(clknet_1_1__leaf_net925),
    .A3(net940),
    .S0(clknet_1_0__leaf_net928),
    .S1(net691),
    .X(net415));
 sky130_fd_sc_hd__a2111o_1 c496 (.A1(net372),
    .A2(clknet_1_0__leaf_net928),
    .B1(clknet_1_0__leaf_net288),
    .C1(clknet_1_1__leaf_net294),
    .D1(net798),
    .X(net416));
 sky130_fd_sc_hd__a2111o_1 c497 (.A1(net409),
    .A2(net978),
    .B1(clknet_1_0__leaf_net288),
    .C1(net875),
    .D1(net695),
    .X(net417));
 sky130_fd_sc_hd__buf_1 c498 (.A(clknet_1_0__leaf_net741),
    .X(net907));
 sky130_fd_sc_hd__and3_1 c499 (.A(net691),
    .B(net892),
    .C(net798),
    .X(net418));
 sky130_fd_sc_hd__a2111o_1 c500 (.A1(clknet_1_1__leaf_net400),
    .A2(clknet_1_0__leaf_net415),
    .B1(clknet_1_0__leaf_net904),
    .C1(net411),
    .D1(net798),
    .X(net419));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net418),
    .A1(net135),
    .A2(net914),
    .A3(net398),
    .S0(net411),
    .S1(net780),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_1__leaf_net151),
    .A1(net420),
    .A2(net411),
    .A3(net398),
    .S0(net691),
    .S1(net780),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(clknet_1_1__leaf_net267),
    .A1(clknet_1_1__leaf_net421),
    .A2(net413),
    .A3(clknet_1_0__leaf_net904),
    .S1(net798),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net135),
    .A1(clknet_1_0__leaf_net421),
    .A2(clknet_1_1__leaf_net288),
    .A3(net923),
    .S0(net420),
    .S1(net757),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_0__leaf_net421),
    .A1(net420),
    .A2(net900),
    .A3(net757),
    .S0(net780),
    .S1(net798),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net985),
    .A1(clknet_1_1__leaf_net264),
    .A2(net885),
    .A3(net940),
    .S0(net71),
    .S1(clknet_1_1__leaf_net925),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net37),
    .A1(net945),
    .A2(net875),
    .A3(clknet_1_1__leaf_net908),
    .S1(net756),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 c528 (.A(net701),
    .X(net427));
 sky130_fd_sc_hd__and2_2 c529 (.A(net209),
    .B(net323),
    .X(net428));
 sky130_fd_sc_hd__buf_1 c530 (.A(net701),
    .X(net429));
 sky130_fd_sc_hd__and2_2 c531 (.A(net195),
    .B(net681),
    .X(net881));
 sky130_fd_sc_hd__dlymetal6s2s_1 c532 (.A(net746),
    .X(net430));
 sky130_fd_sc_hd__and2_1 c533 (.A(net323),
    .B(net332),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 c534 (.A(net700),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c535 (.A(net700),
    .X(net433));
 sky130_fd_sc_hd__a2111o_2 c536 (.A1(net429),
    .A2(net430),
    .B1(net432),
    .C1(net941),
    .D1(net681),
    .X(net434));
 sky130_fd_sc_hd__and2_1 c537 (.A(net427),
    .B(net433),
    .X(net435));
 sky130_fd_sc_hd__and2_4 c538 (.A(net435),
    .B(net433),
    .X(net436));
 sky130_fd_sc_hd__buf_2 c539 (.A(net746),
    .X(net437));
 sky130_fd_sc_hd__sdfbbp_1 c540 (.CLK(clknet_4_1_0_clk),
    .D(net433),
    .RESET_B(net431),
    .SCD(net437),
    .SCE(net432),
    .SET_B(net1009),
    .Q(net439),
    .Q_N(net438));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net195),
    .A1(net439),
    .A2(net437),
    .A3(net431),
    .S0(net209),
    .S1(net881),
    .X(net440));
 sky130_fd_sc_hd__and3_2 c542 (.A(net439),
    .B(net437),
    .C(net792),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net324),
    .A1(net436),
    .A2(net441),
    .A3(net432),
    .S0(net434),
    .S1(net438),
    .X(net442));
 sky130_fd_sc_hd__and2_1 c544 (.A(net439),
    .B(net777),
    .X(net443));
 sky130_fd_sc_hd__a2111o_4 c545 (.A1(net443),
    .A2(net441),
    .B1(net429),
    .C1(net82),
    .D1(net777),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net435),
    .A1(net429),
    .A2(net208),
    .A3(net444),
    .S0(net428),
    .S1(net436),
    .X(net445));
 sky130_fd_sc_hd__a2111o_1 c547 (.A1(net208),
    .A2(net196),
    .B1(net432),
    .C1(net438),
    .D1(net800),
    .X(net446));
 sky130_fd_sc_hd__mux4_2 c548 (.A0(net434),
    .A1(net438),
    .A2(net432),
    .A3(net444),
    .S0(net437),
    .S1(net998),
    .X(net447));
 sky130_fd_sc_hd__mux4_2 c549 (.A0(net446),
    .A1(net84),
    .A2(net444),
    .A3(net447),
    .S0(net441),
    .S1(net800),
    .X(net448));
 sky130_fd_sc_hd__a2111o_4 c550 (.A1(net965),
    .A2(net942),
    .B1(net444),
    .C1(net447),
    .D1(net792),
    .X(net449));
 sky130_fd_sc_hd__or4bb_1 c551 (.A(net942),
    .B(net224),
    .C_N(net965),
    .D_N(net941),
    .X(net450));
 sky130_fd_sc_hd__and3_1 c552 (.A(net82),
    .B(net199),
    .C(net791),
    .X(net451));
 sky130_fd_sc_hd__and2_1 c553 (.A(net427),
    .B(net444),
    .X(net452));
 sky130_fd_sc_hd__and3_4 c554 (.A(net84),
    .B(net953),
    .C(net800),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 c555 (.A(net713),
    .X(net453));
 sky130_fd_sc_hd__buf_1 c556 (.A(net713),
    .X(net454));
 sky130_fd_sc_hd__a2111o_1 c557 (.A1(net446),
    .A2(net941),
    .B1(net449),
    .C1(net956),
    .D1(net905),
    .X(net455));
 sky130_fd_sc_hd__and2_0 c558 (.A(net449),
    .B(net453),
    .X(net456));
 sky130_fd_sc_hd__and3_1 c559 (.A(net453),
    .B(net456),
    .C(net85),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net347),
    .A1(net350),
    .A2(net942),
    .A3(net449),
    .S0(net791),
    .S1(net998),
    .X(net458));
 sky130_fd_sc_hd__and2_1 c561 (.A(net456),
    .B(net821),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net349),
    .A1(net342),
    .A2(net942),
    .A3(net449),
    .S0(net821),
    .S1(net800),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 c563 (.A(net713),
    .X(net461));
 sky130_fd_sc_hd__buf_1 c564 (.A(net713),
    .X(net891));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net450),
    .A1(net350),
    .A2(net459),
    .A3(net948),
    .S0(net446),
    .S1(net949),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net439),
    .A1(net457),
    .A2(net452),
    .A3(net436),
    .S0(net905),
    .S1(net801),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(net455),
    .A1(net447),
    .A2(net463),
    .A3(net448),
    .S0(net347),
    .S1(net801),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net456),
    .A1(net460),
    .A2(net453),
    .A3(net457),
    .S0(net719),
    .S1(net801),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net457),
    .A1(net949),
    .A2(net948),
    .A3(net449),
    .S0(net224),
    .S1(net696),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net463),
    .A1(net454),
    .A2(net448),
    .A3(net235),
    .S0(net778),
    .S1(net801),
    .X(net467));
 sky130_fd_sc_hd__a2111o_2 c571 (.A1(net455),
    .A2(net950),
    .B1(net905),
    .C1(net696),
    .D1(net801),
    .X(net468));
 sky130_fd_sc_hd__and2_0 c572 (.A(net357),
    .B(net828),
    .X(net469));
 sky130_fd_sc_hd__or4bb_4 c573 (.A(net890),
    .B(net949),
    .C_N(net952),
    .D_N(net919),
    .X(net470));
 sky130_fd_sc_hd__and2_0 c574 (.A(net469),
    .B(net199),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net366),
    .A1(net243),
    .A2(net451),
    .A3(net342),
    .S0(net949),
    .S1(net963),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net776),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 c577 (.A(net725),
    .X(net474));
 sky130_fd_sc_hd__and2_0 c578 (.A(net452),
    .B(net1),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net473),
    .A1(net199),
    .A2(net469),
    .A3(net470),
    .S0(net950),
    .S1(net952),
    .X(net476));
 sky130_fd_sc_hd__and2_1 c580 (.A(net474),
    .B(net476),
    .X(net477));
 sky130_fd_sc_hd__and3_1 c581 (.A(net950),
    .B(net379),
    .C(net719),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net451),
    .A1(net477),
    .A2(net430),
    .A3(net478),
    .S0(net468),
    .S1(net357),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net478),
    .A1(net447),
    .A2(net475),
    .A3(net384),
    .S0(net950),
    .S1(net952),
    .X(net480));
 sky130_fd_sc_hd__or4bb_1 c584 (.A(net476),
    .B(net950),
    .C_N(net953),
    .D_N(net919),
    .X(net481));
 sky130_fd_sc_hd__and3_2 c585 (.A(net199),
    .B(net481),
    .C(net357),
    .X(net482));
 sky130_fd_sc_hd__buf_1 c586 (.A(net725),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_1 c587 (.A(net726),
    .X(net483));
 sky130_fd_sc_hd__and2_0 c588 (.A(net481),
    .B(net124),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_2 c589 (.A(net767),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net459),
    .A1(net238),
    .A2(net485),
    .A3(net470),
    .S0(net482),
    .S1(net1),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net483),
    .A1(net870),
    .A2(net485),
    .A3(net477),
    .S0(net482),
    .S1(net1004),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net936),
    .A1(net473),
    .A2(net485),
    .A3(net444),
    .S0(net724),
    .S1(net888),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net947),
    .A1(net485),
    .A2(net905),
    .A3(net724),
    .S0(net888),
    .S1(net801),
    .X(net489));
 sky130_fd_sc_hd__and3_2 c594 (.A(net447),
    .B(net485),
    .C(net828),
    .X(net490));
 sky130_fd_sc_hd__and3_1 c595 (.A(net485),
    .B(net902),
    .C(net755),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 c596 (.A(net897),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 c597 (.A(net897),
    .X(net493));
 sky130_fd_sc_hd__a2111o_1 c598 (.A1(net132),
    .A2(net394),
    .B1(net491),
    .C1(net377),
    .D1(net732),
    .X(net494));
 sky130_fd_sc_hd__buf_1 c599 (.A(net776),
    .X(net893));
 sky130_fd_sc_hd__a2111o_1 c600 (.A1(net475),
    .A2(net490),
    .B1(net491),
    .C1(net905),
    .D1(net132),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c601 (.A(net127),
    .B(net390),
    .C(net491),
    .X(net496));
 sky130_fd_sc_hd__buf_1 c602 (.A(clknet_1_1__leaf_net770),
    .X(net497));
 sky130_fd_sc_hd__a2111o_1 c603 (.A1(net496),
    .A2(net905),
    .B1(net243),
    .C1(clknet_1_1__leaf_net930),
    .D1(net489),
    .X(net498));
 sky130_fd_sc_hd__and3_1 c604 (.A(net370),
    .B(net390),
    .C(net905),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net495),
    .A1(net447),
    .A2(net379),
    .A3(net946),
    .S0(net697),
    .S1(clknet_1_0__leaf_net740),
    .X(net911));
 sky130_fd_sc_hd__and3_1 c606 (.A(net471),
    .B(net71),
    .C(net132),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 c607 (.A(net894),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 c608 (.A(net894),
    .X(net502));
 sky130_fd_sc_hd__and3_1 c609 (.A(net501),
    .B(net946),
    .C(net732),
    .X(net503));
 sky130_fd_sc_hd__a2111o_1 c610 (.A1(net503),
    .A2(net490),
    .B1(net951),
    .C1(net243),
    .D1(net493),
    .X(net504));
 sky130_fd_sc_hd__or4bb_1 c611 (.A(net491),
    .B(net502),
    .C_N(net504),
    .D_N(net951),
    .X(net505));
 sky130_fd_sc_hd__a2111o_1 c612 (.A1(net504),
    .A2(net468),
    .B1(net503),
    .C1(net490),
    .D1(clknet_1_0__leaf_net770),
    .X(net506));
 sky130_fd_sc_hd__a2111o_1 c613 (.A1(net489),
    .A2(net497),
    .B1(net502),
    .C1(net390),
    .D1(net243),
    .X(net507));
 sky130_fd_sc_hd__a2111o_1 c614 (.A1(net390),
    .A2(net470),
    .B1(net732),
    .C1(clknet_1_0__leaf_net770),
    .D1(net776),
    .X(net508));
 sky130_fd_sc_hd__sdfbbn_1 c615 (.CLK_N(clknet_4_3_0_clk),
    .D(net1007),
    .RESET_B(net507),
    .SCD(net492),
    .SCE(net503),
    .SET_B(net490),
    .Q(net510),
    .Q_N(net509));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(clknet_1_0__leaf_net302),
    .A1(net385),
    .A2(net905),
    .A3(net946),
    .S0(net165),
    .S1(net799),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net171),
    .A1(net944),
    .A2(clknet_1_0__leaf_net302),
    .A3(net902),
    .S0(clknet_1_0__leaf_net294),
    .S1(net799),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(clknet_1_0__leaf_net511),
    .A1(net901),
    .A2(net881),
    .A3(net411),
    .S0(net944),
    .S1(net828),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net477),
    .A1(net384),
    .A2(clknet_1_0__leaf_net173),
    .A3(clknet_1_0__leaf_net880),
    .S0(net948),
    .S1(net804),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net868),
    .A1(net873),
    .A2(net876),
    .A3(net962),
    .S0(net864),
    .S1(net869),
    .X(net0));
 sky130_fd_sc_hd__a2111o_1 c620 (.A1(net494),
    .A2(net902),
    .B1(net893),
    .C1(net470),
    .D1(net956),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net413),
    .A1(net499),
    .A2(clknet_1_0__leaf_net907),
    .A3(net420),
    .S0(net951),
    .S1(net804),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net166),
    .A1(clknet_1_1__leaf_net511),
    .A2(net477),
    .A3(net367),
    .S0(clknet_1_1__leaf_net302),
    .S1(net895),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(clknet_1_0__leaf_net151),
    .A1(net468),
    .A2(net74),
    .A3(clknet_1_1__leaf_net508),
    .S0(clknet_1_0__leaf_net908),
    .S1(net899),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(clknet_1_1__leaf_net173),
    .A1(clknet_1_1__leaf_net930),
    .A2(net976),
    .A3(clknet_1_1__leaf_net904),
    .S0(clknet_1_1__leaf_net908),
    .S1(net945),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net367),
    .A1(net411),
    .A2(clknet_1_0__leaf_net511),
    .A3(net470),
    .S0(net420),
    .S1(clknet_1_1__leaf_net512),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net468),
    .A1(clknet_1_0__leaf_net173),
    .A2(net870),
    .A3(clknet_1_0__leaf_net907),
    .S0(net804),
    .S1(net912),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net470),
    .A1(net477),
    .A2(net515),
    .A3(net901),
    .S0(clknet_1_1__leaf_net930),
    .S1(clknet_1_0__leaf_net173),
    .X(net522));
 sky130_fd_sc_hd__a2111o_1 c628 (.A1(net963),
    .A2(net747),
    .B1(net892),
    .C1(net773),
    .D1(net895),
    .X(net523));
 sky130_fd_sc_hd__a2111o_1 c629 (.A1(clknet_1_0__leaf_net294),
    .A2(net875),
    .B1(net948),
    .C1(net515),
    .D1(net912),
    .X(net524));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net860),
    .A1(net862),
    .A2(net869),
    .A3(net0),
    .S0(net849),
    .S1(net961),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net516),
    .A1(net828),
    .A2(net870),
    .A3(clknet_1_1__leaf_net880),
    .S0(net411),
    .S1(net799),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net298),
    .A1(net367),
    .A2(clknet_1_1__leaf_net524),
    .A3(clknet_1_1__leaf_net508),
    .S0(net935),
    .S1(net805),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net875),
    .A1(net509),
    .A2(clknet_1_0__leaf_net908),
    .A3(net926),
    .S0(net895),
    .S1(net805),
    .X(net527));
 sky130_fd_sc_hd__sdfbbn_1 c633 (.CLK_N(clknet_4_8_0_clk),
    .D(clknet_1_1__leaf_net302),
    .RESET_B(clknet_1_1__leaf_net524),
    .SCD(net297),
    .SCE(net894),
    .SET_B(net766),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__a2111o_1 c634 (.A1(net528),
    .A2(clknet_1_1__leaf_net524),
    .B1(net773),
    .C1(net799),
    .D1(net805),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net523),
    .A1(net529),
    .A2(clknet_1_1__leaf_net524),
    .A3(net747),
    .S0(net775),
    .S1(net805),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net528),
    .A1(net436),
    .A2(clknet_1_0__leaf_net930),
    .A3(net695),
    .S0(net736),
    .S1(net775),
    .X(net532));
 sky130_fd_sc_hd__a2111o_1 c637 (.A1(net529),
    .A2(net510),
    .B1(net736),
    .C1(net773),
    .D1(net775),
    .X(net533));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net3),
    .A1(net829),
    .A2(net864),
    .A3(net868),
    .S0(net844),
    .S1(net878),
    .X(net2));
 sky130_fd_sc_hd__mux4_1 c65 (.A0(net878),
    .A1(net835),
    .A2(net842),
    .A3(net845),
    .S0(net843),
    .S1(net829),
    .X(net3));
 sky130_fd_sc_hd__and2_0 c66 (.A(net855),
    .B(net844),
    .X(net4));
 sky130_fd_sc_hd__and2_1 c660 (.A(net443),
    .B(net436),
    .X(net534));
 sky130_fd_sc_hd__and3_1 c661 (.A(net434),
    .B(net441),
    .C(net941),
    .X(net535));
 sky130_fd_sc_hd__buf_1 c662 (.A(net714),
    .X(net536));
 sky130_fd_sc_hd__and2_1 c663 (.A(net536),
    .B(net448),
    .X(net537));
 sky130_fd_sc_hd__and2_0 c664 (.A(net832),
    .B(net535),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_1 c665 (.A(net772),
    .X(net539));
 sky130_fd_sc_hd__and2_0 c666 (.A(net429),
    .B(net535),
    .X(net540));
 sky130_fd_sc_hd__and2_2 c667 (.A(net538),
    .B(net536),
    .X(net541));
 sky130_fd_sc_hd__buf_1 c668 (.A(net772),
    .X(net542));
 sky130_fd_sc_hd__and2_1 c669 (.A(net539),
    .B(net943),
    .X(net543));
 sky130_fd_sc_hd__and2_0 c67 (.A(net824),
    .B(net961),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 c670 (.A(net714),
    .X(net544));
 sky130_fd_sc_hd__or4bb_1 c671 (.A(net540),
    .B(net434),
    .C_N(net542),
    .D_N(net943),
    .X(net545));
 sky130_fd_sc_hd__and2_1 c672 (.A(net432),
    .B(net543),
    .X(net546));
 sky130_fd_sc_hd__and2_0 c673 (.A(net535),
    .B(net546),
    .X(net547));
 sky130_fd_sc_hd__or4bb_4 c674 (.A(net434),
    .B(net939),
    .C_N(net448),
    .D_N(net777),
    .X(net548));
 sky130_fd_sc_hd__or4bb_1 c675 (.A(net545),
    .B(net543),
    .C_N(net548),
    .D_N(net939),
    .X(net549));
 sky130_fd_sc_hd__and3_1 c676 (.A(net535),
    .B(net939),
    .C(net764),
    .X(net550));
 sky130_fd_sc_hd__a2111o_1 c677 (.A1(net543),
    .A2(net542),
    .B1(net546),
    .C1(net939),
    .D1(net832),
    .X(net551));
 sky130_fd_sc_hd__or4bb_1 c678 (.A(net544),
    .B(net536),
    .C_N(net537),
    .D_N(net550),
    .X(net552));
 sky130_fd_sc_hd__a2111o_1 c679 (.A1(net551),
    .A2(net542),
    .B1(net535),
    .C1(net548),
    .X(net553));
 sky130_fd_sc_hd__and2_0 c68 (.A(net2),
    .B(net862),
    .X(net6));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net332),
    .A2(net551),
    .B1(net543),
    .C1(net939),
    .D1(net764),
    .X(net554));
 sky130_fd_sc_hd__sdfbbp_1 c681 (.CLK(clknet_4_0_0_clk),
    .D(net554),
    .RESET_B(net551),
    .SCD(net448),
    .SCE(net536),
    .SET_B(net764),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__a2111o_1 c682 (.A1(net448),
    .A2(net454),
    .B1(net546),
    .C1(net449),
    .D1(net939),
    .X(net557));
 sky130_fd_sc_hd__buf_1 c683 (.A(net727),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net84),
    .A1(net546),
    .A2(net449),
    .A3(net821),
    .S0(net548),
    .S1(net792),
    .X(net559));
 sky130_fd_sc_hd__buf_1 c685 (.A(net727),
    .X(net560));
 sky130_fd_sc_hd__and3_1 c686 (.A(net546),
    .B(net550),
    .C(net448),
    .X(net561));
 sky130_fd_sc_hd__sdfbbn_1 c687 (.CLK_N(clknet_4_1_0_clk),
    .D(net541),
    .RESET_B(net350),
    .SCD(net560),
    .SCE(net683),
    .SET_B(clknet_1_0__leaf_net806),
    .Q(net563),
    .Q_N(net562));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net557),
    .A1(net550),
    .A2(net85),
    .A3(net561),
    .S0(net792),
    .S1(net801),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net548),
    .A1(net556),
    .A2(net560),
    .A3(net546),
    .S0(net937),
    .S1(net449),
    .X(net565));
 sky130_fd_sc_hd__and2_1 c69 (.A(net5),
    .B(net876),
    .X(net7));
 sky130_fd_sc_hd__and3_1 c690 (.A(net941),
    .B(net852),
    .C(net943),
    .X(net566));
 sky130_fd_sc_hd__a2111o_1 c691 (.A1(net550),
    .A2(net828),
    .B1(net556),
    .C1(net941),
    .D1(net954),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net1002),
    .A1(net561),
    .A2(net1012),
    .A3(net550),
    .S0(net937),
    .S1(net801),
    .X(net568));
 sky130_fd_sc_hd__a2111o_1 c693 (.A1(net224),
    .A2(net548),
    .B1(net955),
    .C1(net949),
    .D1(net801),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(net567),
    .A1(net437),
    .A2(net548),
    .A3(net941),
    .S0(net955),
    .S1(net560),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net821),
    .A1(net563),
    .A2(net949),
    .A3(net939),
    .S0(net791),
    .S1(clknet_1_1__leaf_net806),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 c696 (.A(net726),
    .X(net572));
 sky130_fd_sc_hd__and3_1 c697 (.A(net551),
    .B(net778),
    .C(clknet_1_0__leaf_net807),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net573),
    .A1(clknet_1_0__leaf_net571),
    .A2(net554),
    .A3(net550),
    .S0(net572),
    .S1(net792),
    .X(net574));
 sky130_fd_sc_hd__and3_1 c699 (.A(net561),
    .B(net778),
    .C(clknet_1_0__leaf_net808),
    .X(net575));
 sky130_fd_sc_hd__and2_0 c70 (.A(net849),
    .B(net851),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net350),
    .A1(net466),
    .A2(net572),
    .A3(net949),
    .S0(clknet_1_0__leaf_net806),
    .S1(net810),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net561),
    .A1(net554),
    .A2(net555),
    .A3(net714),
    .S0(clknet_1_0__leaf_net808),
    .S1(net812),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net449),
    .A1(net556),
    .A2(clknet_1_0__leaf_net571),
    .A3(net941),
    .S0(net745),
    .S1(clknet_1_0__leaf_net807),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net578),
    .A1(net558),
    .A2(net557),
    .A3(net714),
    .S0(net812),
    .S1(net813),
    .X(net579));
 sky130_fd_sc_hd__or4bb_2 c704 (.A(net563),
    .B(net852),
    .C_N(net541),
    .D_N(net955),
    .X(net580));
 sky130_fd_sc_hd__or4bb_1 c705 (.A(net943),
    .B(net945),
    .C_N(net801),
    .D_N(clknet_1_0__leaf_net808),
    .X(net581));
 sky130_fd_sc_hd__or4bb_1 c706 (.A(net1),
    .B(net581),
    .C_N(net949),
    .D_N(net803),
    .X(net582));
 sky130_fd_sc_hd__buf_2 c707 (.A(net723),
    .X(net583));
 sky130_fd_sc_hd__a2111o_1 c708 (.A1(net583),
    .A2(net943),
    .B1(clknet_1_0__leaf_net582),
    .C1(clknet_1_1__leaf_net807),
    .D1(net811),
    .X(net584));
 sky130_fd_sc_hd__and3_1 c709 (.A(net558),
    .B(net947),
    .C(net541),
    .X(net585));
 sky130_fd_sc_hd__and2_0 c71 (.A(net8),
    .B(net861),
    .X(net9));
 sky130_fd_sc_hd__and3_1 c710 (.A(net430),
    .B(net583),
    .C(net779),
    .X(net586));
 sky130_fd_sc_hd__or4bb_1 c711 (.A(net466),
    .B(net585),
    .C_N(net938),
    .D_N(net1010),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net566),
    .A1(clknet_1_0__leaf_net582),
    .A2(net938),
    .A3(net746),
    .S0(clknet_1_1__leaf_net807),
    .S1(clknet_1_0__leaf_net808),
    .X(net588));
 sky130_fd_sc_hd__or4bb_1 c713 (.A(net351),
    .B(net943),
    .C_N(net558),
    .D_N(net586),
    .X(net589));
 sky130_fd_sc_hd__mux4_2 c714 (.A0(net541),
    .A1(net583),
    .A2(net585),
    .A3(net955),
    .S0(net938),
    .S1(net745),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net85),
    .A1(net945),
    .A2(net437),
    .A3(net590),
    .S0(net947),
    .S1(clknet_1_1__leaf_net807),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_1__leaf_net571),
    .A1(net948),
    .A2(net938),
    .A3(net572),
    .S0(net583),
    .S1(net949),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net590),
    .A1(net558),
    .A2(net541),
    .A3(net572),
    .S0(net803),
    .S1(net815),
    .X(net593));
 sky130_fd_sc_hd__buf_1 c718 (.A(net723),
    .X(net933));
 sky130_fd_sc_hd__and3_1 c719 (.A(net437),
    .B(net592),
    .C(net124),
    .X(net594));
 sky130_fd_sc_hd__and2_2 c72 (.A(net842),
    .B(net874),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net943),
    .A1(net586),
    .A2(net558),
    .A3(net933),
    .S0(net562),
    .S1(net815),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net594),
    .A1(net590),
    .A2(net436),
    .A3(net943),
    .S0(net727),
    .S1(net814),
    .X(net596));
 sky130_fd_sc_hd__a2111o_1 c722 (.A1(net595),
    .A2(net380),
    .B1(net943),
    .C1(net815),
    .D1(net816),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net454),
    .A1(net590),
    .A2(net534),
    .A3(net852),
    .S0(net814),
    .S1(net815),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net588),
    .A1(net590),
    .A2(net937),
    .A3(clknet_1_0__leaf_net582),
    .S0(net1004),
    .S1(net816),
    .X(net599));
 sky130_fd_sc_hd__a2111o_1 c725 (.A1(net597),
    .A2(net727),
    .B1(net771),
    .C1(net809),
    .D1(net816),
    .X(net600));
 sky130_fd_sc_hd__sdfbbn_1 c726 (.CLK_N(clknet_4_2_0_clk),
    .D(net585),
    .RESET_B(net938),
    .SCD(net937),
    .SCE(net852),
    .SET_B(net1001),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__a2111o_1 c727 (.A1(net956),
    .A2(net947),
    .B1(net948),
    .C1(net938),
    .D1(net755),
    .X(net603));
 sky130_fd_sc_hd__or4bb_1 c728 (.A(net938),
    .B(net600),
    .C_N(net585),
    .D_N(net811),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net395),
    .A1(net951),
    .A2(clknet_1_1__leaf_net582),
    .A3(net938),
    .S0(net947),
    .S1(clknet_1_1__leaf_net808),
    .X(net605));
 sky130_fd_sc_hd__and2_0 c73 (.A(net851),
    .B(net6),
    .X(net11));
 sky130_fd_sc_hd__or4bb_1 c730 (.A(net390),
    .B(net124),
    .C_N(net779),
    .D_N(clknet_1_1__leaf_net808),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net601),
    .A1(net503),
    .A2(clknet_1_0__leaf_net508),
    .A3(net937),
    .S0(net938),
    .S1(net743),
    .X(net607));
 sky130_fd_sc_hd__sdfsbp_2 c732 (.CLK(clknet_4_2_0_clk),
    .D(net585),
    .SCD(net937),
    .SCE(net947),
    .SET_B(net817),
    .Q(net609),
    .Q_N(net608));
 sky130_fd_sc_hd__or4bb_1 c733 (.A(net947),
    .B(clknet_1_0__leaf_net584),
    .C_N(net771),
    .D_N(net779),
    .X(net610));
 sky130_fd_sc_hd__or4bb_1 c734 (.A(net955),
    .B(net603),
    .C_N(net608),
    .D_N(clknet_1_1__leaf_net808),
    .X(net611));
 sky130_fd_sc_hd__sdfbbp_1 c735 (.CLK(clknet_4_3_0_clk),
    .D(net380),
    .RESET_B(net238),
    .SCD(clknet_1_1__leaf_net508),
    .SCE(net1008),
    .SET_B(net996),
    .Q(net613),
    .Q_N(net612));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net613),
    .A1(clknet_1_0__leaf_net611),
    .A2(net379),
    .A3(net938),
    .S0(clknet_1_0__leaf_net610),
    .S1(net812),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net613),
    .A1(net609),
    .A2(clknet_1_0__leaf_net614),
    .A3(net379),
    .S0(net746),
    .S1(net810),
    .X(net615));
 sky130_fd_sc_hd__a2111o_1 c738 (.A1(net124),
    .A2(net947),
    .B1(net583),
    .C1(net603),
    .D1(net813),
    .X(net616));
 sky130_fd_sc_hd__a2111o_1 c739 (.A1(net606),
    .A2(net379),
    .B1(net608),
    .C1(net715),
    .D1(net750),
    .X(net617));
 sky130_fd_sc_hd__and2_0 c74 (.A(net11),
    .B(net10),
    .X(net12));
 sky130_fd_sc_hd__a2111o_1 c740 (.A1(net604),
    .A2(clknet_1_1__leaf_net584),
    .B1(clknet_1_0__leaf_net611),
    .C1(net612),
    .D1(net743),
    .X(net618));
 sky130_fd_sc_hd__or4bb_1 c741 (.A(net617),
    .B(clknet_1_1__leaf_net614),
    .C_N(net609),
    .D_N(net750),
    .X(net619));
 sky130_fd_sc_hd__a2111o_1 c742 (.A1(clknet_1_1__leaf_net611),
    .A2(net500),
    .B1(net613),
    .C1(net380),
    .D1(net509),
    .X(net620));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(net238),
    .A2(net616),
    .B1(net956),
    .C1(clknet_1_1__leaf_net611),
    .D1(net814),
    .X(net621));
 sky130_fd_sc_hd__mux4_2 c744 (.A0(net937),
    .A1(net1011),
    .A2(net997),
    .A3(net948),
    .S0(net715),
    .S1(net753),
    .X(net622));
 sky130_fd_sc_hd__or4bb_1 c745 (.A(net616),
    .B(clknet_1_0__leaf_net614),
    .C_N(net753),
    .D_N(net777),
    .X(net623));
 sky130_fd_sc_hd__a2111o_1 c746 (.A1(clknet_1_1__leaf_net610),
    .A2(net608),
    .B1(net600),
    .C1(net716),
    .D1(net777),
    .X(net624));
 sky130_fd_sc_hd__a2111o_1 c747 (.A1(net620),
    .A2(clknet_1_0__leaf_net624),
    .B1(net939),
    .C1(net890),
    .D1(net777),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(clknet_1_1__leaf_net614),
    .A1(net609),
    .A2(clknet_1_0__leaf_net930),
    .A3(net955),
    .S0(net883),
    .S1(net817),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_1__leaf_net605),
    .A1(net533),
    .A2(net436),
    .A3(net744),
    .S0(net799),
    .S1(net935),
    .X(net627));
 sky130_fd_sc_hd__and2_2 c75 (.A(net0),
    .B(net5),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(clknet_1_0__leaf_net508),
    .A1(net890),
    .A2(net609),
    .A3(net947),
    .S0(net951),
    .S1(net817),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net603),
    .A1(net602),
    .A2(clknet_1_0__leaf_net930),
    .A3(clknet_1_0__leaf_net508),
    .S0(net436),
    .S1(net817),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_0__leaf_net605),
    .A1(clknet_1_0__leaf_net628),
    .A2(net602),
    .A3(clknet_1_0__leaf_net880),
    .S0(clknet_1_0__leaf_net508),
    .S1(net951),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_0__leaf_net512),
    .A1(net490),
    .A2(clknet_1_1__leaf_net582),
    .A3(net934),
    .S0(net979),
    .S1(net935),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net946),
    .A1(net852),
    .A2(net948),
    .A3(clknet_1_0__leaf_net624),
    .S0(clknet_1_0__leaf_net930),
    .S1(net816),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net948),
    .A1(net881),
    .A2(net934),
    .A3(net411),
    .S0(net963),
    .S1(net888),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(clknet_1_0__leaf_net524),
    .A1(net627),
    .A2(net74),
    .A3(clknet_1_0__leaf_net508),
    .S0(net775),
    .S1(net817),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net436),
    .A1(net533),
    .A2(net609),
    .A3(net515),
    .S0(clknet_1_0__leaf_net508),
    .S1(net580),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net493),
    .A1(net411),
    .A2(net603),
    .A3(net890),
    .S0(net980),
    .S1(net818),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net583),
    .A1(clknet_1_0__leaf_net151),
    .A2(clknet_1_0__leaf_net880),
    .A3(clknet_1_0__leaf_net524),
    .S0(net744),
    .S1(net900),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c76 (.A0(net8),
    .A1(net859),
    .A2(net13),
    .A3(net10),
    .S0(net826),
    .S1(net872),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net515),
    .A1(net71),
    .A2(net420),
    .A3(clknet_1_1__leaf_net624),
    .S0(net377),
    .S1(clknet_1_0__leaf_net512),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(clknet_1_0__leaf_net151),
    .A1(net946),
    .A2(clknet_1_1__leaf_net508),
    .A3(clknet_1_0__leaf_net930),
    .S0(net533),
    .S1(net818),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(clknet_1_1__leaf_net582),
    .A1(net934),
    .A2(clknet_1_0__leaf_net880),
    .A3(net891),
    .S0(net892),
    .S1(net766),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net636),
    .A1(net635),
    .A2(clknet_1_0__leaf_net524),
    .A3(net963),
    .S0(net601),
    .S1(clknet_1_1__leaf_net628),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net420),
    .A1(net411),
    .A2(net951),
    .A3(clknet_1_1__leaf_net582),
    .S0(net608),
    .S1(net775),
    .X(net882));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(clknet_1_1__leaf_net624),
    .A1(net749),
    .A2(net919),
    .A3(net883),
    .S0(net799),
    .S1(net818),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net385),
    .A1(net633),
    .A2(net932),
    .A3(clknet_1_1__leaf_net642),
    .S0(net944),
    .S1(net818),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net951),
    .A1(clknet_1_1__leaf_net642),
    .A2(clknet_1_1__leaf_net643),
    .A3(net510),
    .S0(clknet_1_0__leaf_net930),
    .S1(net816),
    .X(net644));
 sky130_fd_sc_hd__a2111o_1 c768 (.A1(net580),
    .A2(clknet_1_0__leaf_net642),
    .B1(clknet_1_0__leaf_net643),
    .C1(net749),
    .D1(net775),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net510),
    .A1(clknet_1_0__leaf_net643),
    .A2(net645),
    .A3(clknet_1_0__leaf_net642),
    .S0(net956),
    .S1(net716),
    .X(net646));
 sky130_fd_sc_hd__and2_2 c77 (.A(net14),
    .B(net874),
    .X(net910));
 sky130_fd_sc_hd__and2_1 c78 (.A(net874),
    .B(net861),
    .X(net15));
 sky130_fd_sc_hd__and2_0 c79 (.A(net9),
    .B(net962),
    .X(net16));
 sky130_fd_sc_hd__and3_2 c80 (.A(net13),
    .B(net14),
    .C(net861),
    .X(net17));
 sky130_fd_sc_hd__and3_1 c81 (.A(net16),
    .B(net858),
    .C(net2),
    .X(net18));
 sky130_fd_sc_hd__and3_1 c82 (.A(net857),
    .B(net18),
    .C(net14),
    .X(net19));
 sky130_fd_sc_hd__or4bb_2 c83 (.A(net12),
    .B(net9),
    .C_N(net10),
    .D_N(net17),
    .X(net20));
 sky130_fd_sc_hd__or4bb_1 c84 (.A(net18),
    .B(net17),
    .C_N(net20),
    .D_N(net7),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net19),
    .A1(net860),
    .A2(net4),
    .A3(net20),
    .S0(net867),
    .S1(net21),
    .X(net22));
 sky130_fd_sc_hd__and3_1 c86 (.A(net17),
    .B(net21),
    .C(net20),
    .X(net23));
 sky130_fd_sc_hd__and3_1 c87 (.A(net21),
    .B(net23),
    .C(net20),
    .X(net24));
 sky130_fd_sc_hd__and2_2 c88 (.A(net867),
    .B(net910),
    .X(net25));
 sky130_fd_sc_hd__and3_1 c89 (.A(net876),
    .B(net25),
    .C(net2),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c90 (.A(net6),
    .B(net946),
    .X(net27));
 sky130_fd_sc_hd__and3_4 c91 (.A(net862),
    .B(net17),
    .C(net23),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c92 (.A(net865),
    .B(net28),
    .X(net29));
 sky130_fd_sc_hd__and2_0 c93 (.A(net23),
    .B(net859),
    .X(net30));
 sky130_fd_sc_hd__and2_4 c94 (.A(net22),
    .B(net25),
    .X(net31));
 sky130_fd_sc_hd__and3_1 c95 (.A(net30),
    .B(net31),
    .C(net27),
    .X(net32));
 sky130_fd_sc_hd__and2_1 c96 (.A(net27),
    .B(net29),
    .X(net33));
 sky130_fd_sc_hd__and2_1 c97 (.A(net32),
    .B(net33),
    .X(net34));
 sky130_fd_sc_hd__and2_1 c98 (.A(net29),
    .B(net34),
    .X(net35));
 sky130_fd_sc_hd__and3_1 c99 (.A(net4),
    .B(net2),
    .C(net865),
    .X(net36));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net406),
    .A1(net367),
    .A2(clknet_1_0__leaf_net264),
    .A3(net134),
    .S0(net969),
    .S1(clknet_1_1__leaf_net768),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net167),
    .A1(clknet_1_1__leaf_net916),
    .A2(clknet_1_1__leaf_net179),
    .A3(net59),
    .S0(net190),
    .S1(net186),
    .X(net648));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net108),
    .A1(net236),
    .A2(net271),
    .A3(net116),
    .S0(net993),
    .S1(net782),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net320),
    .A1(net324),
    .A2(net327),
    .A3(net331),
    .S0(net334),
    .S1(net791),
    .X(net650));
 sky130_fd_sc_hd__or4bb_1 merge794 (.A(net431),
    .B(net535),
    .C_N(net542),
    .D_N(net537),
    .X(net651));
 sky130_fd_sc_hd__mux4_2 merge795 (.A0(net428),
    .A1(net490),
    .A2(net963),
    .A3(net116),
    .S0(net482),
    .S1(net949),
    .X(net652));
 sky130_fd_sc_hd__or4bb_1 merge796 (.A(net342),
    .B(net351),
    .C_N(net936),
    .D_N(net470),
    .X(net653));
 sky130_fd_sc_hd__or4bb_1 merge797 (.A(net320),
    .B(net339),
    .C_N(net327),
    .D_N(net85),
    .X(net654));
 sky130_fd_sc_hd__or4bb_1 merge798 (.A(net235),
    .B(net447),
    .C_N(net234),
    .D_N(net449),
    .X(net655));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net239),
    .A1(net236),
    .A2(net109),
    .A3(net115),
    .S0(net238),
    .S1(net228),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net572),
    .A1(net466),
    .A2(net541),
    .A3(net590),
    .S0(net562),
    .S1(net1003),
    .X(net657));
 sky130_fd_sc_hd__a2111o_1 merge801 (.A1(clknet_1_0__leaf_net284),
    .A2(net922),
    .B1(clknet_1_1__leaf_net880),
    .C1(net291),
    .D1(net923),
    .X(net658));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net939),
    .A1(net557),
    .A2(net554),
    .A3(net937),
    .S0(net555),
    .S1(net791),
    .X(net659));
 sky130_fd_sc_hd__or4bb_1 merge803 (.A(net55),
    .B(net2),
    .C_N(net845),
    .D_N(net57),
    .X(net660));
 sky130_fd_sc_hd__a2111o_1 merge804 (.A1(net836),
    .A2(net10),
    .B1(net984),
    .C1(net139),
    .D1(net24),
    .X(net661));
 sky130_fd_sc_hd__or4bb_1 merge805 (.A(net428),
    .B(net427),
    .C_N(net825),
    .D_N(net339),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge806 (.A0(net1021),
    .A1(net973),
    .A2(net983),
    .A3(net43),
    .S0(net35),
    .S1(net40),
    .X(net663));
 sky130_fd_sc_hd__a2111o_1 merge807 (.A1(net128),
    .A2(net326),
    .B1(net125),
    .C1(net109),
    .D1(clknet_1_0__leaf_net740),
    .X(net664));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net190),
    .A1(clknet_1_1__leaf_net415),
    .A2(clknet_1_1__leaf_net904),
    .A3(clknet_1_1__leaf_net267),
    .S0(net759),
    .S1(net788),
    .X(net665));
 sky130_fd_sc_hd__or4bb_1 merge809 (.A(net221),
    .B(net226),
    .C_N(net343),
    .D_N(net953),
    .X(net666));
 sky130_fd_sc_hd__a2111o_1 merge810 (.A1(net480),
    .A2(net482),
    .B1(net561),
    .C1(net821),
    .D1(net809),
    .X(net667));
 sky130_fd_sc_hd__a2111o_1 merge811 (.A1(net472),
    .A2(net492),
    .B1(net490),
    .C1(net444),
    .D1(net238),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 merge812 (.A0(net472),
    .A1(clknet_1_0__leaf_net277),
    .A2(net270),
    .A3(net386),
    .S0(net697),
    .S1(net732),
    .X(net669));
 sky130_fd_sc_hd__a2111o_1 merge813 (.A1(net339),
    .A2(net431),
    .B1(net77),
    .C1(net332),
    .D1(net428),
    .X(net670));
 sky130_fd_sc_hd__a2111o_1 merge814 (.A1(net450),
    .A2(net890),
    .B1(net954),
    .C1(net460),
    .D1(net459),
    .X(net671));
 sky130_fd_sc_hd__a2111o_1 merge815 (.A1(net537),
    .A2(net332),
    .B1(net943),
    .C1(net441),
    .D1(net832),
    .X(net672));
 sky130_fd_sc_hd__mux4_1 merge816 (.A0(net109),
    .A1(net351),
    .A2(net936),
    .A3(net482),
    .S0(net946),
    .S1(net963),
    .X(net673));
 sky130_fd_sc_hd__mux4_1 merge817 (.A0(net247),
    .A1(net245),
    .A2(net249),
    .A3(net484),
    .S0(net366),
    .S1(net936),
    .X(net674));
 sky130_fd_sc_hd__and2_0 merge818 (.A(net549),
    .B(net552),
    .X(net675));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net615),
    .B(net618),
    .X(net676));
 sky130_fd_sc_hd__and2_0 merge820 (.A(net514),
    .B(net517),
    .X(net677));
 sky130_fd_sc_hd__and2_0 merge821 (.A(net646),
    .B(net626),
    .X(net678));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net61),
    .B(net65),
    .X(net679));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net479),
    .B(net488),
    .X(net680));
 sky130_fd_sc_hd__dfrbp_1 merge824 (.CLK(clknet_4_4_0_clk),
    .D(net325),
    .RESET_B(net336),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dfrbp_1 merge825 (.CLK(clknet_4_5_0_clk),
    .D(net346),
    .RESET_B(net355),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__and2_0 merge826 (.A(net498),
    .B(net505),
    .X(net685));
 sky130_fd_sc_hd__and2_0 merge827 (.A(net257),
    .B(net258),
    .X(net686));
 sky130_fd_sc_hd__dfrtn_1 merge828 (.CLK_N(clknet_4_7_0_clk),
    .D(net666),
    .RESET_B(net233),
    .Q(net687));
 sky130_fd_sc_hd__and2_0 merge829 (.A(net569),
    .B(net574),
    .X(net688));
 sky130_fd_sc_hd__and2_0 merge830 (.A(net140),
    .B(net142),
    .X(net689));
 sky130_fd_sc_hd__and2_0 merge831 (.A(net155),
    .B(net168),
    .X(net690));
 sky130_fd_sc_hd__dfrtp_4 merge832 (.CLK(clknet_4_15_0_clk),
    .D(net45),
    .RESET_B(net42),
    .Q(net691));
 sky130_fd_sc_hd__and2_0 merge833 (.A(net387),
    .B(net404),
    .X(net692));
 sky130_fd_sc_hd__and2_0 merge834 (.A(net295),
    .B(net299),
    .X(net693));
 sky130_fd_sc_hd__and2_0 merge835 (.A(net305),
    .B(net306),
    .X(net694));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_4_11_0_clk),
    .D(net425),
    .Q(net426));
 sky130_fd_sc_hd__dfrtp_1 merge837 (.CLK(clknet_4_9_0_clk),
    .D(net412),
    .RESET_B(net410),
    .Q(net695));
 sky130_fd_sc_hd__dfsbp_1 merge838 (.CLK(clknet_4_1_0_clk),
    .D(net464),
    .SET_B(net465),
    .Q(net697),
    .Q_N(net696));
 sky130_fd_sc_hd__and2_0 merge839 (.A(net213),
    .B(net212),
    .X(net698));
 sky130_fd_sc_hd__and2_0 merge840 (.A(net587),
    .B(net598),
    .X(net699));
 sky130_fd_sc_hd__dfsbp_1 merge841 (.CLK(clknet_4_4_0_clk),
    .D(net654),
    .SET_B(net662),
    .Q(net701),
    .Q_N(net700));
 sky130_fd_sc_hd__and2_0 merge842 (.A(net269),
    .B(net273),
    .X(net702));
 sky130_fd_sc_hd__and2_0 merge843 (.A(net192),
    .B(net194),
    .X(net703));
 sky130_fd_sc_hd__and2_0 merge844 (.A(net378),
    .B(net382),
    .X(net704));
 sky130_fd_sc_hd__and2_0 merge845 (.A(net527),
    .B(net518),
    .X(net705));
 sky130_fd_sc_hd__and2_0 merge846 (.A(net278),
    .B(net405),
    .X(net706));
 sky130_fd_sc_hd__and2_0 merge847 (.A(net634),
    .B(net678),
    .X(net707));
 sky130_fd_sc_hd__and2_0 merge848 (.A(net506),
    .B(net673),
    .X(net708));
 sky130_fd_sc_hd__dfstp_1 merge849 (.CLK(clknet_4_5_0_clk),
    .D(net664),
    .SET_B(net650),
    .Q(net709));
 sky130_fd_sc_hd__and2_0 merge850 (.A(net621),
    .B(net638),
    .X(net710));
 sky130_fd_sc_hd__and2_0 merge851 (.A(net575),
    .B(net579),
    .X(net711));
 sky130_fd_sc_hd__and2_0 merge852 (.A(net644),
    .B(net641),
    .X(net712));
 sky130_fd_sc_hd__dfstp_1 merge853 (.CLK(clknet_4_4_0_clk),
    .D(net671),
    .SET_B(net655),
    .Q(net713));
 sky130_fd_sc_hd__dfstp_1 merge854 (.CLK(clknet_4_0_0_clk),
    .D(net651),
    .SET_B(net688),
    .Q(net714));
 sky130_fd_sc_hd__dlrbn_1 merge855 (.D(net710),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net676),
    .Q(net716),
    .Q_N(net715));
 sky130_fd_sc_hd__and2_0 merge856 (.A(net150),
    .B(net702),
    .X(net717));
 sky130_fd_sc_hd__dlrbn_1 merge857 (.D(net359),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net352),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__and2_0 merge858 (.A(net313),
    .B(net308),
    .X(net720));
 sky130_fd_sc_hd__and2_0 merge859 (.A(net316),
    .B(net522),
    .X(net721));
 sky130_fd_sc_hd__and2_0 merge860 (.A(net526),
    .B(net639),
    .X(net722));
 sky130_fd_sc_hd__dlrbp_1 merge861 (.D(net680),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net657),
    .Q(net724),
    .Q_N(net723));
 sky130_fd_sc_hd__dlrbp_1 merge862 (.D(net667),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net653),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__dlrtn_1 merge863 (.D(net659),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net699),
    .Q(net727));
 sky130_fd_sc_hd__and2_0 merge864 (.A(net629),
    .B(net632),
    .X(net728));
 sky130_fd_sc_hd__and2_0 merge865 (.A(net137),
    .B(net661),
    .X(net729));
 sky130_fd_sc_hd__dlrtn_2 merge866 (.D(net728),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net487),
    .Q(net888));
 sky130_fd_sc_hd__and2_0 merge867 (.A(net312),
    .B(net174),
    .X(net730));
 sky130_fd_sc_hd__and2_0 merge868 (.A(net656),
    .B(net674),
    .X(net731));
 sky130_fd_sc_hd__dlrtn_2 merge869 (.D(net698),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net232),
    .Q(net732));
 sky130_fd_sc_hd__and2_0 merge870 (.A(net309),
    .B(net317),
    .X(net733));
 sky130_fd_sc_hd__dlrtp_1 merge871 (.D(net663),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net690),
    .Q(net734));
 sky130_fd_sc_hd__dlrtp_1 merge872 (.GATE(clknet_4_6_0_clk),
    .RESET_B(net704),
    .Q(net381));
 sky130_fd_sc_hd__dlrtp_1 merge873 (.D(net310),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net531),
    .Q(net736));
 sky130_fd_sc_hd__edfxbp_1 merge874 (.CLK(clknet_4_12_0_clk),
    .D(net692),
    .DE(net706),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__edfxtp_1 merge875 (.CLK(clknet_4_15_0_clk),
    .D(net184),
    .DE(net733),
    .Q(net739));
 sky130_fd_sc_hd__sdlclkp_1 merge876 (.CLK(clknet_4_7_0_clk),
    .GATE(net689),
    .SCE(net126),
    .GCLK(net740));
 sky130_fd_sc_hd__sdlclkp_2 merge877 (.CLK(clknet_4_11_0_clk),
    .GATE(net703),
    .SCE(net665),
    .GCLK(net741));
 sky130_fd_sc_hd__sdlclkp_4 merge878 (.CLK(clknet_4_12_0_clk),
    .GATE(net268),
    .SCE(net658),
    .GCLK(net742));
 sky130_fd_sc_hd__dfrbp_1 merge879 (.CLK(clknet_4_8_0_clk),
    .D(net593),
    .RESET_B(net721),
    .Q(net743),
    .Q_N(net926));
 sky130_fd_sc_hd__dfrbp_1 merge880 (.CLK(clknet_4_2_0_clk),
    .D(net711),
    .RESET_B(net625),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dfrtn_1 merge881 (.CLK_N(clknet_4_0_0_clk),
    .D(net670),
    .RESET_B(net568),
    .Q(net746));
 sky130_fd_sc_hd__dfrtp_2 merge882 (.CLK(clknet_4_12_0_clk),
    .D(net293),
    .RESET_B(net414),
    .Q(net747));
 sky130_fd_sc_hd__dfrtp_1 merge883 (.CLK(clknet_4_14_0_clk),
    .D(net189),
    .RESET_B(net283),
    .Q(net748));
 sky130_fd_sc_hd__dfrtp_4 merge884 (.CLK(clknet_4_13_0_clk),
    .D(net652),
    .RESET_B(net730),
    .Q(net897));
 sky130_fd_sc_hd__dfsbp_1 merge885 (.CLK(clknet_4_2_0_clk),
    .D(net589),
    .SET_B(net712),
    .Q(net750),
    .Q_N(net749));
 sky130_fd_sc_hd__dfsbp_1 merge886 (.CLK(clknet_4_14_0_clk),
    .D(net693),
    .SET_B(net720),
    .Q(net751),
    .Q_N(net886));
 sky130_fd_sc_hd__dfstp_1 merge887 (.CLK(clknet_4_10_0_clk),
    .D(net423),
    .SET_B(net707),
    .Q(net900));
 sky130_fd_sc_hd__dfstp_1 merge888 (.CLK(clknet_4_12_0_clk),
    .D(net647),
    .SET_B(net649),
    .Q(net752));
 sky130_fd_sc_hd__dfstp_2 merge889 (.CLK(clknet_4_3_0_clk),
    .D(net467),
    .SET_B(net623),
    .Q(net919));
 sky130_fd_sc_hd__dlrbn_1 merge890 (.D(net619),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net694),
    .Q(net753),
    .Q_N(net921));
 sky130_fd_sc_hd__dlrbn_1 merge891 (.D(net261),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net686),
    .Q(net755),
    .Q_N(net754));
 sky130_fd_sc_hd__dlrbp_1 merge892 (.GATE(clknet_4_11_0_clk),
    .RESET_B(net417),
    .Q(net757),
    .Q_N(net756));
 sky130_fd_sc_hd__dlrbp_1 merge893 (.D(net181),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net648),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__and2_0 merge894 (.A(net315),
    .B(net187),
    .X(net760));
 sky130_fd_sc_hd__dlrtn_1 merge895 (.D(net668),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net705),
    .Q(net894));
 sky130_fd_sc_hd__dlrtn_1 merge896 (.D(net307),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net660),
    .Q(net761));
 sky130_fd_sc_hd__dlrtn_2 merge897 (.D(net353),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net375),
    .Q(net762));
 sky130_fd_sc_hd__dlrtp_2 merge898 (.D(net637),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net416),
    .Q(net892));
 sky130_fd_sc_hd__dlrtp_2 merge899 (.D(net356),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net358),
    .Q(net763));
 sky130_fd_sc_hd__dlrtp_1 merge900 (.GATE(clknet_4_0_0_clk),
    .RESET_B(net675),
    .Q(net553));
 sky130_fd_sc_hd__and2_0 merge901 (.A(net640),
    .B(net631),
    .X(net765));
 sky130_fd_sc_hd__edfxbp_1 merge902 (.CLK(clknet_4_10_0_clk),
    .D(net722),
    .DE(net677),
    .Q(net766),
    .Q_N(net899));
 sky130_fd_sc_hd__edfxtp_1 merge903 (.CLK(clknet_4_7_0_clk),
    .D(net256),
    .DE(net731),
    .Q(net767));
 sky130_fd_sc_hd__sdlclkp_1 merge904 (.CLK(clknet_4_12_0_clk),
    .GATE(net717),
    .SCE(net403),
    .GCLK(net768));
 sky130_fd_sc_hd__sdlclkp_2 merge905 (.CLK(clknet_4_15_0_clk),
    .GATE(net679),
    .SCE(net276),
    .GCLK(net769));
 sky130_fd_sc_hd__sdlclkp_4 merge906 (.CLK(clknet_4_9_0_clk),
    .GATE(net685),
    .SCE(net669),
    .GCLK(net770));
 sky130_fd_sc_hd__dfrbp_1 merge907 (.CLK(clknet_4_3_0_clk),
    .D(net672),
    .RESET_B(net599),
    .Q(net772),
    .Q_N(net771));
 sky130_fd_sc_hd__dfrbp_2 merge908 (.CLK(clknet_4_10_0_clk),
    .D(net521),
    .RESET_B(net532),
    .Q(net773),
    .Q_N(net883));
 sky130_fd_sc_hd__dfrtn_1 merge909 (.CLK_N(clknet_4_13_0_clk),
    .D(net279),
    .RESET_B(net729),
    .Q(net774));
 sky130_fd_sc_hd__dfrtp_4 merge910 (.CLK(clknet_4_10_0_clk),
    .D(net765),
    .RESET_B(net530),
    .Q(net775));
 sky130_fd_sc_hd__dfrtp_4 merge911 (.CLK(clknet_4_11_0_clk),
    .D(net708),
    .RESET_B(net760),
    .Q(net776));
 sky130_fd_sc_hd__dfrtp_4 merge912 (.CLK(clknet_4_1_0_clk),
    .D(net442),
    .RESET_B(net622),
    .Q(net777));
 sky130_fd_sc_hd__dfsbp_1 merge913 (.CLK(clknet_4_1_0_clk),
    .D(net440),
    .SET_B(net458),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__dfsbp_1 merge914 (.CLK(clknet_4_11_0_clk),
    .D(net60),
    .SET_B(net419),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dfxbp_1 s915 (.CLK(clknet_4_13_0_clk),
    .D(net147),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_4_13_0_clk),
    .D(net148),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dfxtp_1 s917 (.CLK(clknet_4_13_0_clk),
    .D(net149),
    .Q(net786));
 sky130_fd_sc_hd__dfxtp_1 s918 (.CLK(clknet_4_15_0_clk),
    .D(net183),
    .Q(net787));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_4_15_0_clk),
    .D(net188),
    .Q(net788));
 sky130_fd_sc_hd__dlclkp_1 s920 (.CLK(clknet_4_7_0_clk),
    .GATE(net250),
    .GCLK(net789));
 sky130_fd_sc_hd__dlclkp_2 s921 (.CLK(clknet_4_7_0_clk),
    .GATE(net254),
    .GCLK(net790));
 sky130_fd_sc_hd__dlclkp_4 s922 (.CLK(clknet_4_14_0_clk),
    .GATE(net296),
    .GCLK(net931));
 sky130_fd_sc_hd__dlxbn_2 s923 (.D(net333),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net337),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net794),
    .Q_N(net793));
 sky130_fd_sc_hd__dlxbp_1 s925 (.D(net383),
    .GATE(clknet_4_6_0_clk),
    .Q(net796),
    .Q_N(net795));
 sky130_fd_sc_hd__dlxtn_1 s926 (.D(net402),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net797));
 sky130_fd_sc_hd__dlxtn_2 s927 (.D(net407),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net798));
 sky130_fd_sc_hd__dlxtn_2 s928 (.D(net424),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net799));
 sky130_fd_sc_hd__dlxtp_1 s929 (.D(net445),
    .GATE(clknet_4_4_0_clk),
    .Q(net800));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s930 (.D(net462),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net801));
 sky130_fd_sc_hd__dfxbp_1 s931 (.CLK(clknet_4_3_0_clk),
    .D(net486),
    .Q(net803),
    .Q_N(net802));
 sky130_fd_sc_hd__dfxbp_1 s932 (.CLK(clknet_4_9_0_clk),
    .D(net513),
    .Q(net895),
    .Q_N(net804));
 sky130_fd_sc_hd__dfxtp_2 s933 (.CLK(clknet_4_11_0_clk),
    .D(net519),
    .Q(net935));
 sky130_fd_sc_hd__dfxtp_1 s934 (.CLK(clknet_4_9_0_clk),
    .D(net520),
    .Q(net912));
 sky130_fd_sc_hd__dfxtp_1 s935 (.CLK(clknet_4_10_0_clk),
    .D(net525),
    .Q(net805));
 sky130_fd_sc_hd__dlclkp_1 s936 (.CLK(clknet_4_1_0_clk),
    .GATE(net559),
    .GCLK(net806));
 sky130_fd_sc_hd__dlclkp_2 s937 (.CLK(clknet_4_0_0_clk),
    .GATE(net564),
    .GCLK(net807));
 sky130_fd_sc_hd__dlclkp_4 s938 (.CLK(clknet_4_0_0_clk),
    .GATE(net565),
    .GCLK(net808));
 sky130_fd_sc_hd__dlxbn_1 s939 (.D(net570),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dlxbn_1 s940 (.D(net576),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net812),
    .Q_N(net811));
 sky130_fd_sc_hd__dlxbp_1 s941 (.D(net577),
    .GATE(clknet_4_0_0_clk),
    .Q(net814),
    .Q_N(net813));
 sky130_fd_sc_hd__dlxtn_1 s942 (.D(net591),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net815));
 sky130_fd_sc_hd__dlxtn_2 s943 (.D(net596),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net816));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net607),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net817));
 sky130_fd_sc_hd__dlxtp_1 s945 (.D(net630),
    .GATE(clknet_4_8_0_clk),
    .Q(net818));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net422));
 sky130_fd_sc_hd__buf_6 input2 (.A(in1),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net821));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(in12),
    .X(net822));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(in13),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net824));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net827));
 sky130_fd_sc_hd__buf_4 input11 (.A(in18),
    .X(net828));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input14 (.A(in20),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in22),
    .X(net833));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net834));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in25),
    .X(net836));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input24 (.A(in3),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net842));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net843));
 sky130_fd_sc_hd__buf_2 input27 (.A(in32),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net845));
 sky130_fd_sc_hd__buf_6 input29 (.A(in34),
    .X(net846));
 sky130_fd_sc_hd__buf_6 input30 (.A(in35),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in36),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net851));
 sky130_fd_sc_hd__buf_4 input35 (.A(in4),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in40),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net854));
 sky130_fd_sc_hd__buf_2 input38 (.A(in42),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net856));
 sky130_fd_sc_hd__buf_1 input40 (.A(in44),
    .X(net857));
 sky130_fd_sc_hd__buf_2 input41 (.A(in45),
    .X(net858));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input47 (.A(in50),
    .X(net864));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(in51),
    .X(net865));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net866));
 sky130_fd_sc_hd__buf_1 input50 (.A(in53),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net868));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(in56),
    .X(net870));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net871));
 sky130_fd_sc_hd__buf_2 input55 (.A(in58),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net873));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net874));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net875));
 sky130_fd_sc_hd__buf_1 input59 (.A(in61),
    .X(net876));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net877));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(in8),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in9),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(clknet_1_0__leaf_net880),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output64 (.A(net881),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net882),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net883),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net884),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output68 (.A(net885),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net886),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net955),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net888),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net981),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net890),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output74 (.A(net948),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net892),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output76 (.A(net893),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net894),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output78 (.A(net895),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output79 (.A(net974),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output80 (.A(net897),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(clknet_1_1__leaf_net898),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output82 (.A(net899),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output83 (.A(net900),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output84 (.A(net901),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output85 (.A(net902),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output86 (.A(net903),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(clknet_1_1__leaf_net904),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output88 (.A(net905),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output89 (.A(net906),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(clknet_1_1__leaf_net907),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(clknet_1_1__leaf_net908),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output92 (.A(net909),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net910),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net911),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output95 (.A(net912),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net913),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output97 (.A(net914),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output98 (.A(net915),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(clknet_1_0__leaf_net916),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output100 (.A(net917),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output101 (.A(net918),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output102 (.A(net919),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net920),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output104 (.A(net921),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output105 (.A(net940),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output106 (.A(net923),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(clknet_1_1__leaf_net924),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(clknet_1_1__leaf_net925),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output109 (.A(net926),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net927),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(clknet_1_1__leaf_net928),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net929),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(clknet_1_0__leaf_net930),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net931),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output115 (.A(net932),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output116 (.A(net933),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output117 (.A(net947),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output118 (.A(net935),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(net371),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net231),
    .X(net937));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net547),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net922),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net203),
    .X(net941));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net318),
    .X(net942));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(net534),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net910),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net906),
    .X(net945));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net7),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net934),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net891),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net951),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net461),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net732),
    .X(net952));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net341),
    .X(net954));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net887),
    .X(net955));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net887),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net960),
    .X(net957));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_8 fanout142 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(net87),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net867),
    .X(net961));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net866),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net855),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net808 (.A(net808),
    .X(clknet_0_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_0__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_1__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net614 (.A(net614),
    .X(clknet_0_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_0__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net614 (.A(clknet_0_net614),
    .X(clknet_1_1__leaf_net614));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net582 (.A(net582),
    .X(clknet_0_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_0__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_1__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net610 (.A(net610),
    .X(clknet_0_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_0__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net610 (.A(clknet_0_net610),
    .X(clknet_1_1__leaf_net610));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net624 (.A(net624),
    .X(clknet_0_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net624 (.A(clknet_0_net624),
    .X(clknet_1_0__leaf_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net624 (.A(clknet_0_net624),
    .X(clknet_1_1__leaf_net624));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net642 (.A(net642),
    .X(clknet_0_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_0__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net642 (.A(clknet_0_net642),
    .X(clknet_1_1__leaf_net642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net643 (.A(net643),
    .X(clknet_0_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_0__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net643 (.A(clknet_0_net643),
    .X(clknet_1_1__leaf_net643));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net807 (.A(net807),
    .X(clknet_0_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_0__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net807 (.A(clknet_0_net807),
    .X(clknet_1_1__leaf_net807));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net806 (.A(net806),
    .X(clknet_0_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_0__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_1__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net512 (.A(net512),
    .X(clknet_0_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_0__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net512 (.A(clknet_0_net512),
    .X(clknet_1_1__leaf_net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net511 (.A(net511),
    .X(clknet_0_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_0__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net511 (.A(clknet_0_net511),
    .X(clknet_1_1__leaf_net511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net790 (.A(net790),
    .X(clknet_0_net790));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net790 (.A(clknet_0_net790),
    .X(clknet_1_0__leaf_net790));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net790 (.A(clknet_0_net790),
    .X(clknet_1_1__leaf_net790));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net789 (.A(net789),
    .X(clknet_0_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_0__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_1__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net741 (.A(net741),
    .X(clknet_0_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_0__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net741 (.A(clknet_0_net741),
    .X(clknet_1_1__leaf_net741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net907 (.A(net907),
    .X(clknet_0_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_0__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net907 (.A(clknet_0_net907),
    .X(clknet_1_1__leaf_net907));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net908 (.A(net908),
    .X(clknet_0_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_1__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net277 (.A(net277),
    .X(clknet_0_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_0__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net277 (.A(clknet_0_net277),
    .X(clknet_1_1__leaf_net277));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net770 (.A(net770),
    .X(clknet_0_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_1__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net508 (.A(net508),
    .X(clknet_0_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_0__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net508 (.A(clknet_0_net508),
    .X(clknet_1_1__leaf_net508));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net628 (.A(net628),
    .X(clknet_0_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_0__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net628 (.A(clknet_0_net628),
    .X(clknet_1_1__leaf_net628));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net930 (.A(net930),
    .X(clknet_0_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net524 (.A(net524),
    .X(clknet_0_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_0__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net524 (.A(clknet_0_net524),
    .X(clknet_1_1__leaf_net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net263 (.A(net263),
    .X(clknet_0_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_0__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net263 (.A(clknet_0_net263),
    .X(clknet_1_1__leaf_net263));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net285 (.A(net285),
    .X(clknet_0_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_0__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net285 (.A(clknet_0_net285),
    .X(clknet_1_1__leaf_net285));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net288 (.A(net288),
    .X(clknet_0_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_0__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net288 (.A(clknet_0_net288),
    .X(clknet_1_1__leaf_net288));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net284 (.A(net284),
    .X(clknet_0_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_0__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net284 (.A(clknet_0_net284),
    .X(clknet_1_1__leaf_net284));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net768 (.A(net768),
    .X(clknet_0_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_0__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net768 (.A(clknet_0_net768),
    .X(clknet_1_1__leaf_net768));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net275 (.A(net275),
    .X(clknet_0_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_0__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net275 (.A(clknet_0_net275),
    .X(clknet_1_1__leaf_net275));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net63 (.A(net63),
    .X(clknet_0_net63));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net63 (.A(clknet_0_net63),
    .X(clknet_1_0__leaf_net63));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net63 (.A(clknet_0_net63),
    .X(clknet_1_1__leaf_net63));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net267 (.A(net267),
    .X(clknet_0_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net267 (.A(clknet_0_net267),
    .X(clknet_1_0__leaf_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net267 (.A(net982),
    .X(clknet_1_1__leaf_net267));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net928 (.A(net928),
    .X(clknet_0_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net928 (.A(clknet_0_net928),
    .X(clknet_1_0__leaf_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net928 (.A(clknet_0_net928),
    .X(clknet_1_1__leaf_net928));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net415 (.A(net415),
    .X(clknet_0_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_0__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_1__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net400 (.A(net400),
    .X(clknet_0_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_0__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net400 (.A(clknet_0_net400),
    .X(clknet_1_1__leaf_net400));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net252 (.A(net252),
    .X(clknet_0_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_0__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net252 (.A(clknet_0_net252),
    .X(clknet_1_1__leaf_net252));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net253 (.A(net253),
    .X(clknet_0_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_0__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_1__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net264 (.A(net264),
    .X(clknet_0_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_0__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net264 (.A(clknet_0_net264),
    .X(clknet_1_1__leaf_net264));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net740 (.A(net740),
    .X(clknet_0_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_0__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net740 (.A(clknet_0_net740),
    .X(clknet_1_1__leaf_net740));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net916 (.A(net916),
    .X(clknet_0_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_0__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_1__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net913 (.A(net913),
    .X(clknet_0_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_0__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net913 (.A(clknet_0_net913),
    .X(clknet_1_1__leaf_net913));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net152 (.A(net152),
    .X(clknet_0_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_0__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_1__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net281 (.A(net281),
    .X(clknet_0_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_0__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net281 (.A(clknet_0_net281),
    .X(clknet_1_1__leaf_net281));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net880 (.A(net880),
    .X(clknet_0_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net173 (.A(net173),
    .X(clknet_0_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_0__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net173 (.A(clknet_0_net173),
    .X(clknet_1_1__leaf_net173));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net151 (.A(net151),
    .X(clknet_0_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_0__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net151 (.A(clknet_0_net151),
    .X(clknet_1_1__leaf_net151));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net104),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net964),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net112),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net966),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net98),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net1018),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net87),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net896),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net896),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net972),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net972),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net974),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net974),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net972),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net889),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net978),
    .X(net979));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer17 (.A(net979),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net889),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(clknet_0_net267),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net134),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net983),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_1 clone22 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net87),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net960),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net987),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(net959),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_1 clone27 (.A(net960),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(clknet_1_0__leaf_net267),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net991),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(net992),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net734),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net763),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net772),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net612),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net800),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net365),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net762),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net810),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net560),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net811),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net802),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net292),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net792),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net374),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net394),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net435),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net803),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net395),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net437),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net763),
    .X(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_D_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_B (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_D_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_C1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_D_N (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_SCD (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_D1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_C_N (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_RESET_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_D (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_RESET_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S0 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_SCD (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_X (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_Q_N (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_Q (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_D_N (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_D_N (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_C (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_C (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_C1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_RESET_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_D_N (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_D (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_RESET_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_D1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_D1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_C1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_SCE (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_C_N (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_D1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_SET_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_X (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_C1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_D (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_RESET_B (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_C1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_X (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_Q_N (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_C1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_D (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_Q (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_Q_N (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_C1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_Q (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_C1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_B1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_X (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_D1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S0 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCD (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_X (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_C1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_D_N (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A0 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_C1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_X (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_D_N (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_C1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_D (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_RESET_B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_X (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_B1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_X (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_RESET_B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_X (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_D (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_X (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_RESET_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_Q (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_SET_B (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_C (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_Q (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D_N (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_SET_B (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_C (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_RESET_B (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_X (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_D1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_C (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_S1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_Q (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_B1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_D_N (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCD (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_Q (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_Q (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_C1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_Q (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_C (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_D_N (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_D1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_D1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_Q (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_C_N (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_Q (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_D1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_D1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_D_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_Q (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCE (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_C (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D_N (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge910_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_D1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_D1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_Q (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_D1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_D1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_C_N (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_Q (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_D1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_D1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_D_N (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_D_N (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_D1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_Q (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_D_N (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_C_N (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_C (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_C1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_D_N (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_C (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_Q (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_D1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_C (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_C1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_C (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_C (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_C_N (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C_N (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_D1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_D1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_D1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_D1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_D1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_D_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_C1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_C (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_C (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_D1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_D1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_D_N (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_C_N (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_C (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_C_N (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCE (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_C (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_C (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_B1 (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_C (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C_N (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_C1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_C1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net880_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge908_Q_N (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_Q (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_C1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_B1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_Q (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_B1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_B1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_Q (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_D1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_Q (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_C (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_Q (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_C (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_C (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_C1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_D1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_D1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_D_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_C_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_Q (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_D_N (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D_N (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_Q_N (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_D_N (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_D1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_RESET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_RESET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_D_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_Q_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_Q (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_Q (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_S1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SCD (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SET_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_C_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCD (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SCE (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_SCD (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_SCD (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_C1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_RESET_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_C_N (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_B1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_D1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_C1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_C1 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_D_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_D_N (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_C (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_D_N (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_C (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_D_N (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_C_N (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_RESET_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_D1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_B1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_D_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_C (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_D_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_D_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_D1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SET_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_D_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_C1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_C (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_B1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_D1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_D1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D_N (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_B1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_D1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_C1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_D1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_C (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_SCE (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_SCE (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_SCE (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge900_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge899_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge903_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_D1 (.DIODE(clknet_1_0__leaf_net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(clknet_1_0__leaf_net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D1 (.DIODE(clknet_1_0__leaf_net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net790_X (.DIODE(clknet_1_0__leaf_net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S0 (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net930_X (.DIODE(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A0 (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_C1 (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net930_X (.DIODE(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net880_X (.DIODE(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_B1 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_B1 (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net880_X (.DIODE(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_C1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_C_N (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_RESET_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_C_N (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C_N (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net987));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net107),
    .A1(net104),
    .A2(net92),
    .A3(net83),
    .S0(net1021),
    .S1(net101),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net134),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net134),
    .X(net1016));
 sky130_fd_sc_hd__or4bb_1 clone28 (.A(net97),
    .B(net846),
    .C_N(net839),
    .D_N(net959),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net87),
    .X(net1018));
 sky130_fd_sc_hd__and3_1 clone32 (.A(net819),
    .B(net846),
    .C(net847),
    .X(net1019));
 sky130_fd_sc_hd__and3_1 clone33 (.A(net958),
    .B(net89),
    .C(net854),
    .X(net1020));
 sky130_fd_sc_hd__and3_1 clone34 (.A(net958),
    .B(net89),
    .C(net854),
    .X(net1021));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
