module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net628;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net794;
 wire clknet_1_0__leaf_net794;
 wire clknet_1_1__leaf_net794;
 wire clknet_0_net568;
 wire clknet_1_0__leaf_net568;
 wire clknet_1_1__leaf_net568;
 wire clknet_0_net774;
 wire clknet_1_0__leaf_net774;
 wire clknet_1_1__leaf_net774;
 wire clknet_0_net591;
 wire clknet_1_0__leaf_net591;
 wire clknet_1_1__leaf_net591;
 wire clknet_0_net698;
 wire clknet_1_0__leaf_net698;
 wire clknet_1_1__leaf_net698;
 wire clknet_0_net590;
 wire clknet_1_0__leaf_net590;
 wire clknet_1_1__leaf_net590;
 wire clknet_0_net775;
 wire clknet_1_0__leaf_net775;
 wire clknet_1_1__leaf_net775;
 wire clknet_0_net587;
 wire clknet_1_0__leaf_net587;
 wire clknet_1_1__leaf_net587;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net333;
 wire clknet_1_0__leaf_net333;
 wire clknet_1_1__leaf_net333;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net737;
 wire clknet_1_0__leaf_net737;
 wire clknet_1_1__leaf_net737;
 wire clknet_0_net793;
 wire clknet_1_0__leaf_net793;
 wire clknet_1_1__leaf_net793;
 wire clknet_0_net360;
 wire clknet_1_0__leaf_net360;
 wire clknet_1_1__leaf_net360;
 wire clknet_0_net792;
 wire clknet_1_0__leaf_net792;
 wire clknet_1_1__leaf_net792;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net773;
 wire clknet_1_0__leaf_net773;
 wire clknet_1_1__leaf_net773;
 wire clknet_0_net583;
 wire clknet_1_0__leaf_net583;
 wire clknet_1_1__leaf_net583;
 wire clknet_0_net561;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_1__leaf_net561;
 wire clknet_0_net541;
 wire clknet_1_0__leaf_net541;
 wire clknet_1_1__leaf_net541;
 wire clknet_0_net757;
 wire clknet_1_0__leaf_net757;
 wire clknet_1_1__leaf_net757;
 wire clknet_0_net517;
 wire clknet_1_0__leaf_net517;
 wire clknet_1_1__leaf_net517;
 wire clknet_0_net621;
 wire clknet_1_0__leaf_net621;
 wire clknet_1_1__leaf_net621;
 wire clknet_0_net756;
 wire clknet_1_0__leaf_net756;
 wire clknet_1_1__leaf_net756;
 wire clknet_0_net755;
 wire clknet_1_0__leaf_net755;
 wire clknet_1_1__leaf_net755;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net736;
 wire clknet_1_0__leaf_net736;
 wire clknet_1_1__leaf_net736;
 wire clknet_0_net925;
 wire clknet_1_0__leaf_net925;
 wire clknet_1_1__leaf_net925;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net265;
 wire clknet_1_0__leaf_net265;
 wire clknet_1_1__leaf_net265;
 wire clknet_0_net909;
 wire clknet_1_0__leaf_net909;
 wire clknet_1_1__leaf_net909;
 wire clknet_0_net238;
 wire clknet_1_0__leaf_net238;
 wire clknet_1_1__leaf_net238;
 wire clknet_0_net246;
 wire clknet_1_0__leaf_net246;
 wire clknet_1_1__leaf_net246;
 wire clknet_0_net718;
 wire clknet_1_0__leaf_net718;
 wire clknet_1_1__leaf_net718;
 wire clknet_0_net206;
 wire clknet_1_0__leaf_net206;
 wire clknet_1_1__leaf_net206;
 wire clknet_0_net312;
 wire clknet_1_0__leaf_net312;
 wire clknet_1_1__leaf_net312;
 wire clknet_0_net322;
 wire clknet_1_0__leaf_net322;
 wire clknet_1_1__leaf_net322;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net870;
 wire clknet_1_0__leaf_net870;
 wire clknet_1_1__leaf_net870;
 wire clknet_0_net309;
 wire clknet_1_0__leaf_net309;
 wire clknet_1_1__leaf_net309;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net305;
 wire clknet_1_0__leaf_net305;
 wire clknet_1_1__leaf_net305;
 wire clknet_0_net717;
 wire clknet_1_0__leaf_net717;
 wire clknet_1_1__leaf_net717;
 wire clknet_0_net274;
 wire clknet_1_0__leaf_net274;
 wire clknet_1_1__leaf_net274;
 wire clknet_0_net699;
 wire clknet_1_0__leaf_net699;
 wire clknet_1_1__leaf_net699;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;

 sky130_fd_sc_hd__and2_1 c100 (.A(net31),
    .B(net875),
    .X(net35));
 sky130_fd_sc_hd__and2_2 c101 (.A(net29),
    .B(net11),
    .X(net36));
 sky130_fd_sc_hd__and3_1 c102 (.A(net16),
    .B(net33),
    .C(net31),
    .X(net37));
 sky130_fd_sc_hd__and2_2 c103 (.A(net23),
    .B(net875),
    .X(net910));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net29),
    .A1(net25),
    .A2(net28),
    .A3(net875),
    .S0(net851),
    .S1(net836),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c105 (.A0(net32),
    .A1(net38),
    .A2(net25),
    .A3(net33),
    .S0(net875),
    .S1(net34),
    .X(net888));
 sky130_fd_sc_hd__mux4_2 c106 (.A0(net22),
    .A1(net910),
    .A2(net31),
    .A3(net11),
    .S0(net888),
    .S1(net26),
    .X(net39));
 sky130_fd_sc_hd__and2_0 c107 (.A(net39),
    .B(net38),
    .X(net40));
 sky130_fd_sc_hd__and2_4 c108 (.A(net39),
    .B(net37),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net40),
    .A1(net38),
    .A2(net28),
    .A3(net910),
    .S0(net3),
    .S1(net23),
    .X(net42));
 sky130_fd_sc_hd__and2_0 c110 (.A(net861),
    .B(net851),
    .X(net43));
 sky130_fd_sc_hd__and2_0 c111 (.A(net39),
    .B(net851),
    .X(net44));
 sky130_fd_sc_hd__and2_0 c112 (.A(net958),
    .B(net44),
    .X(net45));
 sky130_fd_sc_hd__and2_1 c113 (.A(net821),
    .B(net34),
    .X(net46));
 sky130_fd_sc_hd__and2_0 c114 (.A(net46),
    .B(net958),
    .X(net47));
 sky130_fd_sc_hd__and2_0 c115 (.A(net25),
    .B(net958),
    .X(net48));
 sky130_fd_sc_hd__and2_1 c116 (.A(net951),
    .B(net47),
    .X(net924));
 sky130_fd_sc_hd__and2_1 c117 (.A(net44),
    .B(net816),
    .X(net49));
 sky130_fd_sc_hd__and2_1 c118 (.A(net31),
    .B(net34),
    .X(net50));
 sky130_fd_sc_hd__and2_1 c119 (.A(net924),
    .B(net50),
    .X(net51));
 sky130_fd_sc_hd__and3_1 c120 (.A(net34),
    .B(net51),
    .C(net49),
    .X(net913));
 sky130_fd_sc_hd__and2_2 c121 (.A(net24),
    .B(net924),
    .X(net52));
 sky130_fd_sc_hd__a2111o_1 c122 (.A1(net49),
    .A2(net50),
    .B1(net31),
    .C1(net851),
    .D1(net52),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c123 (.A(net47),
    .B(net24),
    .X(net54));
 sky130_fd_sc_hd__and2_2 c124 (.A(net43),
    .B(net46),
    .X(net894));
 sky130_fd_sc_hd__and2_0 c125 (.A(net48),
    .B(net49),
    .X(net55));
 sky130_fd_sc_hd__and2_0 c126 (.A(net54),
    .B(net962),
    .X(net56));
 sky130_fd_sc_hd__and2_0 c127 (.A(net53),
    .B(net52),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net57),
    .A1(net53),
    .A2(net52),
    .A3(net55),
    .S0(net894),
    .S1(net49),
    .X(net58));
 sky130_fd_sc_hd__and2_0 c129 (.A(net53),
    .B(net964),
    .X(net904));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net55),
    .A1(net46),
    .A2(net904),
    .A3(net894),
    .S0(net53),
    .X(net59));
 sky130_fd_sc_hd__and2_0 c131 (.A(net56),
    .B(net871),
    .X(net60));
 sky130_fd_sc_hd__and2_1 c132 (.A(net863),
    .B(net813),
    .X(net61));
 sky130_fd_sc_hd__and2_1 c133 (.A(net864),
    .B(net628),
    .X(net62));
 sky130_fd_sc_hd__and2_0 c134 (.A(net61),
    .B(net808),
    .X(net63));
 sky130_fd_sc_hd__and2_2 c135 (.A(net811),
    .B(net61),
    .X(net64));
 sky130_fd_sc_hd__and3_1 c136 (.A(net63),
    .B(net818),
    .C(net809),
    .X(net65));
 sky130_fd_sc_hd__and3_2 c137 (.A(net810),
    .B(net815),
    .C(net863),
    .X(net66));
 sky130_fd_sc_hd__and2_4 c138 (.A(net62),
    .B(net64),
    .X(net67));
 sky130_fd_sc_hd__and2_1 c139 (.A(net628),
    .B(net806),
    .X(net68));
 sky130_fd_sc_hd__and2_1 c140 (.A(net65),
    .B(net814),
    .X(net69));
 sky130_fd_sc_hd__and2_2 c141 (.A(net68),
    .B(net66),
    .X(net70));
 sky130_fd_sc_hd__or4bb_1 c142 (.A(net809),
    .B(net812),
    .C_N(net69),
    .D_N(net817),
    .X(net71));
 sky130_fd_sc_hd__and2_1 c143 (.A(net71),
    .B(net69),
    .X(net72));
 sky130_fd_sc_hd__and2_0 c144 (.A(net827),
    .B(net71),
    .X(net73));
 sky130_fd_sc_hd__or4bb_1 c145 (.A(net72),
    .B(net813),
    .C_N(net68),
    .D_N(net949),
    .X(net74));
 sky130_fd_sc_hd__and2_2 c146 (.A(net69),
    .B(net73),
    .X(net75));
 sky130_fd_sc_hd__and3_1 c147 (.A(net812),
    .B(net64),
    .C(net67),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 c148 (.A0(net66),
    .A1(net76),
    .A2(net65),
    .A3(net827),
    .S0(net864),
    .S1(net67),
    .X(net77));
 sky130_fd_sc_hd__and2_0 c149 (.A(net75),
    .B(net77),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c150 (.A(net77),
    .B(net78),
    .C(net71),
    .X(net79));
 sky130_fd_sc_hd__or4bb_4 c151 (.A(net78),
    .B(net71),
    .C_N(net64),
    .D_N(net812),
    .X(net80));
 sky130_fd_sc_hd__and3_1 c152 (.A(net80),
    .B(net63),
    .C(net76),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net77),
    .A1(net81),
    .A2(net76),
    .A3(net80),
    .S0(net811),
    .S1(net64),
    .X(net869));
 sky130_fd_sc_hd__and2_4 c154 (.A(net819),
    .B(net64),
    .X(net868));
 sky130_fd_sc_hd__and2_2 c155 (.A(net842),
    .B(net68),
    .X(net82));
 sky130_fd_sc_hd__and2_1 c156 (.A(net828),
    .B(net832),
    .X(net83));
 sky130_fd_sc_hd__and2_1 c157 (.A(net73),
    .B(net74),
    .X(net84));
 sky130_fd_sc_hd__and2_0 c158 (.A(net826),
    .B(net82),
    .X(net85));
 sky130_fd_sc_hd__and2_0 c159 (.A(net84),
    .B(net82),
    .X(net86));
 sky130_fd_sc_hd__and2_1 c160 (.A(net85),
    .B(net83),
    .X(net87));
 sky130_fd_sc_hd__and3_2 c161 (.A(net834),
    .B(net868),
    .C(net83),
    .X(net88));
 sky130_fd_sc_hd__and2_1 c162 (.A(net68),
    .B(net805),
    .X(net89));
 sky130_fd_sc_hd__and2_1 c163 (.A(net86),
    .B(net824),
    .X(net90));
 sky130_fd_sc_hd__and3_2 c164 (.A(net807),
    .B(net806),
    .C(net90),
    .X(net91));
 sky130_fd_sc_hd__and3_4 c165 (.A(net841),
    .B(net91),
    .C(net832),
    .X(net92));
 sky130_fd_sc_hd__and2_2 c166 (.A(net63),
    .B(net73),
    .X(net93));
 sky130_fd_sc_hd__and2_2 c167 (.A(net86),
    .B(net92),
    .X(net94));
 sky130_fd_sc_hd__a2111o_1 c168 (.A1(net825),
    .A2(net88),
    .B1(net68),
    .C1(net93),
    .D1(net84),
    .X(net95));
 sky130_fd_sc_hd__a2111o_1 c169 (.A1(net95),
    .A2(net91),
    .B1(net93),
    .C1(net64),
    .D1(net868),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net868),
    .A1(net83),
    .A2(net807),
    .A3(net96),
    .S0(net95),
    .S1(net865),
    .X(net97));
 sky130_fd_sc_hd__and2_1 c171 (.A(net83),
    .B(net91),
    .X(net98));
 sky130_fd_sc_hd__or4bb_1 c172 (.A(net822),
    .B(net85),
    .C_N(net94),
    .D_N(net88),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net97),
    .A1(net69),
    .A2(net82),
    .A3(net92),
    .S0(net94),
    .S1(net91),
    .X(net100));
 sky130_fd_sc_hd__a2111o_4 c174 (.A1(net100),
    .A2(net820),
    .B1(net98),
    .C1(net91),
    .D1(net94),
    .X(net101));
 sky130_fd_sc_hd__sdfbbn_2 c175 (.CLK_N(clknet_4_0_0_clk),
    .D(net833),
    .RESET_B(net100),
    .SCD(net99),
    .SCE(net94),
    .SET_B(net101),
    .Q(net103),
    .Q_N(net102));
 sky130_fd_sc_hd__or4bb_1 c176 (.A(net845),
    .B(net93),
    .C_N(net856),
    .D_N(net3),
    .X(net104));
 sky130_fd_sc_hd__or4bb_2 c177 (.A(net99),
    .B(net858),
    .C_N(net846),
    .D_N(net849),
    .X(net105));
 sky130_fd_sc_hd__buf_1 c178 (.A(net684),
    .X(net106));
 sky130_fd_sc_hd__and3_1 c179 (.A(net859),
    .B(net2),
    .C(net79),
    .X(net107));
 sky130_fd_sc_hd__and3_1 c180 (.A(net107),
    .B(net89),
    .C(net106),
    .X(net108));
 sky130_fd_sc_hd__and3_1 c181 (.A(net69),
    .B(net830),
    .C(net857),
    .X(net109));
 sky130_fd_sc_hd__and3_2 c182 (.A(net0),
    .B(net106),
    .C(net856),
    .X(net110));
 sky130_fd_sc_hd__and3_1 c183 (.A(net830),
    .B(net823),
    .C(net0),
    .X(net111));
 sky130_fd_sc_hd__and3_2 c184 (.A(net846),
    .B(net104),
    .C(net107),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c185 (.A(net106),
    .B(net858),
    .C(net857),
    .X(net113));
 sky130_fd_sc_hd__or4bb_1 c186 (.A(net848),
    .B(net101),
    .C_N(net102),
    .D_N(net940),
    .X(net114));
 sky130_fd_sc_hd__and3_2 c187 (.A(net91),
    .B(net110),
    .C(net940),
    .X(net878));
 sky130_fd_sc_hd__or4bb_4 c188 (.A(net106),
    .B(net110),
    .C_N(net98),
    .D_N(net936),
    .X(net923));
 sky130_fd_sc_hd__and3_1 c189 (.A(net852),
    .B(net936),
    .C(net940),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c190 (.A(net940),
    .B(net805),
    .C(net115),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c191 (.A(net79),
    .B(net94),
    .C(net935),
    .X(net117));
 sky130_fd_sc_hd__or4bb_2 c192 (.A(net116),
    .B(net846),
    .C_N(net110),
    .D_N(net936),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 c193 (.A(net684),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c194 (.A0(net119),
    .A1(net824),
    .A2(net112),
    .A3(net105),
    .S0(net940),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net837),
    .A1(net116),
    .A2(net87),
    .A3(net112),
    .S0(net117),
    .S1(net706),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net104),
    .A1(net116),
    .A2(net121),
    .A3(net119),
    .S0(net67),
    .S1(net940),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net94),
    .A1(net111),
    .A2(net89),
    .A3(net935),
    .S0(net684),
    .S1(net706),
    .X(net123));
 sky130_fd_sc_hd__a2111o_1 c198 (.A1(net1),
    .A2(net918),
    .B1(net856),
    .C1(net121),
    .D1(net108),
    .X(net124));
 sky130_fd_sc_hd__and2_1 c199 (.A(net90),
    .B(net18),
    .X(net125));
 sky130_fd_sc_hd__and3_1 c200 (.A(net823),
    .B(net923),
    .C(net868),
    .X(net126));
 sky130_fd_sc_hd__or4bb_2 c201 (.A(net61),
    .B(net935),
    .C_N(net125),
    .D_N(net940),
    .X(net127));
 sky130_fd_sc_hd__buf_1 c202 (.A(net694),
    .X(net128));
 sky130_fd_sc_hd__and2_1 c203 (.A(net819),
    .B(net19),
    .X(net129));
 sky130_fd_sc_hd__a2111o_2 c204 (.A1(net940),
    .A2(net110),
    .B1(net857),
    .C1(net936),
    .D1(net710),
    .X(net130));
 sky130_fd_sc_hd__or4bb_4 c205 (.A(net129),
    .B(net88),
    .C_N(net130),
    .D_N(net936),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net856),
    .A1(net940),
    .A2(net22),
    .A3(net951),
    .S0(net105),
    .S1(net131),
    .X(net132));
 sky130_fd_sc_hd__or4bb_1 c207 (.A(net849),
    .B(net949),
    .C_N(net812),
    .D_N(net935),
    .X(net133));
 sky130_fd_sc_hd__and2_2 c208 (.A(net133),
    .B(net127),
    .X(net134));
 sky130_fd_sc_hd__a2111o_1 c209 (.A1(net12),
    .A2(net880),
    .B1(net134),
    .C1(net129),
    .D1(net92),
    .X(net135));
 sky130_fd_sc_hd__a2111o_1 c210 (.A1(net13),
    .A2(net940),
    .B1(net923),
    .C1(net960),
    .D1(net92),
    .X(net136));
 sky130_fd_sc_hd__buf_1 c211 (.A(net694),
    .X(net137));
 sky130_fd_sc_hd__or4bb_1 c212 (.A(net959),
    .B(net137),
    .C_N(net850),
    .D_N(net127),
    .X(net138));
 sky130_fd_sc_hd__sdfbbn_1 c213 (.CLK_N(clknet_4_4_0_clk),
    .D(net111),
    .RESET_B(net137),
    .SCD(net138),
    .SCE(net1),
    .SET_B(net135),
    .Q(net140),
    .Q_N(net139));
 sky130_fd_sc_hd__or4bb_4 c214 (.A(net138),
    .B(net108),
    .C_N(net139),
    .D_N(net137),
    .X(net907));
 sky130_fd_sc_hd__a2111o_1 c215 (.A1(net108),
    .A2(net959),
    .B1(net139),
    .C1(net134),
    .D1(net137),
    .X(net141));
 sky130_fd_sc_hd__sdfbbp_1 c216 (.CLK(clknet_4_4_0_clk),
    .D(net135),
    .RESET_B(net141),
    .SCD(net138),
    .SCE(net140),
    .SET_B(net907),
    .Q(net143),
    .Q_N(net142));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(net121),
    .A1(net113),
    .A2(net127),
    .A3(net140),
    .S0(net90),
    .S1(net907),
    .X(net144));
 sky130_fd_sc_hd__a2111o_1 c218 (.A1(net140),
    .A2(net137),
    .B1(net142),
    .C1(net125),
    .D1(net128),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net145),
    .A1(net143),
    .A2(net112),
    .A3(net141),
    .S0(net131),
    .S1(net137),
    .X(net146));
 sky130_fd_sc_hd__and3_1 c220 (.A(net962),
    .B(net27),
    .C(net36),
    .X(net147));
 sky130_fd_sc_hd__or4bb_4 c221 (.A(net18),
    .B(net22),
    .C_N(net142),
    .D_N(net93),
    .X(net898));
 sky130_fd_sc_hd__buf_1 c222 (.A(net996),
    .X(net148));
 sky130_fd_sc_hd__and3_2 c223 (.A(net836),
    .B(net806),
    .C(net898),
    .X(net149));
 sky130_fd_sc_hd__a2111o_1 c224 (.A1(net1),
    .A2(net92),
    .B1(net831),
    .C1(net898),
    .D1(net130),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net898),
    .A1(net851),
    .A2(net843),
    .A3(net134),
    .S0(net42),
    .S1(net706),
    .X(net151));
 sky130_fd_sc_hd__and3_1 c226 (.A(net957),
    .B(net836),
    .C(net26),
    .X(net152));
 sky130_fd_sc_hd__a2111o_4 c227 (.A1(net2),
    .A2(net147),
    .B1(net130),
    .C1(net3),
    .D1(net957),
    .X(net921));
 sky130_fd_sc_hd__and3_2 c228 (.A(net831),
    .B(net143),
    .C(net898),
    .X(net914));
 sky130_fd_sc_hd__and2_0 c229 (.A(net130),
    .B(net147),
    .X(net153));
 sky130_fd_sc_hd__sdfrbp_2 c230 (.CLK(clknet_4_4_0_clk),
    .D(net141),
    .RESET_B(net914),
    .SCD(net149),
    .SCE(net150),
    .Q(net917),
    .Q_N(net154));
 sky130_fd_sc_hd__or4bb_1 c231 (.A(net33),
    .B(net147),
    .C_N(net14),
    .D_N(net152),
    .X(net155));
 sky130_fd_sc_hd__and2_2 c232 (.A(net150),
    .B(net706),
    .X(net156));
 sky130_fd_sc_hd__and2_0 c233 (.A(net152),
    .B(net154),
    .X(net157));
 sky130_fd_sc_hd__buf_1 c234 (.A(net694),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 c235 (.A0(net126),
    .A1(net156),
    .A2(net157),
    .A3(net134),
    .S0(net148),
    .S1(net972),
    .X(net159));
 sky130_fd_sc_hd__sdfbbn_1 c236 (.CLK_N(clknet_4_5_0_clk),
    .D(net156),
    .RESET_B(net158),
    .SCD(net152),
    .SCE(net155),
    .SET_B(net671),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net153),
    .A1(net148),
    .A2(net156),
    .A3(net936),
    .S0(net110),
    .S1(net910),
    .X(net162));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net875),
    .A1(net158),
    .A2(net898),
    .A3(net33),
    .S0(net156),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net148),
    .A1(net910),
    .A2(net2),
    .A3(net1),
    .S0(net156),
    .S1(net126),
    .X(net164));
 sky130_fd_sc_hd__mux4_2 c240 (.A0(net157),
    .A1(net92),
    .A2(net161),
    .A3(net147),
    .S0(net706),
    .S1(net884),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(net165),
    .A1(net152),
    .A2(net151),
    .A3(net671),
    .S0(net715),
    .S1(net884),
    .X(net166));
 sky130_fd_sc_hd__and3_1 c242 (.A(net43),
    .B(net60),
    .C(net49),
    .X(net922));
 sky130_fd_sc_hd__and3_1 c243 (.A(net158),
    .B(net51),
    .C(net914),
    .X(net167));
 sky130_fd_sc_hd__a2111o_1 c244 (.A1(net49),
    .A2(net917),
    .B1(net52),
    .C1(net913),
    .D1(net871),
    .X(net168));
 sky130_fd_sc_hd__and3_1 c245 (.A(net52),
    .B(net894),
    .C(net963),
    .X(net169));
 sky130_fd_sc_hd__or4bb_1 c246 (.A(net806),
    .B(net851),
    .C_N(net907),
    .D_N(net965),
    .X(net170));
 sky130_fd_sc_hd__or4bb_2 c247 (.A(net112),
    .B(net898),
    .C_N(net52),
    .D_N(net715),
    .X(net906));
 sky130_fd_sc_hd__or4bb_2 c248 (.A(net851),
    .B(net93),
    .C_N(net906),
    .D_N(net922),
    .X(net171));
 sky130_fd_sc_hd__and3_1 c249 (.A(net169),
    .B(net910),
    .C(net14),
    .X(net916));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net817),
    .A1(net851),
    .A2(net916),
    .A3(net871),
    .S0(net900),
    .S1(net884),
    .X(net172));
 sky130_fd_sc_hd__and3_1 c251 (.A(net110),
    .B(net910),
    .C(net871),
    .X(net173));
 sky130_fd_sc_hd__and3_2 c252 (.A(net50),
    .B(net906),
    .C(net916),
    .X(net174));
 sky130_fd_sc_hd__a2111o_1 c253 (.A1(net172),
    .A2(net174),
    .B1(net171),
    .C1(net173),
    .D1(net52),
    .X(net175));
 sky130_fd_sc_hd__a2111o_1 c254 (.A1(net173),
    .A2(net966),
    .B1(net907),
    .C1(net174),
    .D1(net997),
    .X(net176));
 sky130_fd_sc_hd__a2111o_2 c255 (.A1(net45),
    .A2(net93),
    .B1(net174),
    .C1(net52),
    .D1(net906),
    .X(net911));
 sky130_fd_sc_hd__and3_1 c256 (.A(net155),
    .B(net174),
    .C(net93),
    .X(net177));
 sky130_fd_sc_hd__sdfrbp_1 c257 (.CLK(clknet_4_5_0_clk),
    .D(net174),
    .RESET_B(net171),
    .SCD(net173),
    .SCE(net900),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net147),
    .A1(net911),
    .A2(net52),
    .A3(net954),
    .S0(net918),
    .S1(net808),
    .X(net905));
 sky130_fd_sc_hd__sdfbbn_1 c259 (.CLK_N(clknet_4_5_0_clk),
    .D(net177),
    .RESET_B(net171),
    .SCD(net911),
    .SCE(net178),
    .SET_B(net154),
    .Q(net181),
    .Q_N(net180));
 sky130_fd_sc_hd__a2111o_1 c260 (.A1(net983),
    .A2(net181),
    .B1(net894),
    .C1(net174),
    .D1(net171),
    .X(net182));
 sky130_fd_sc_hd__a2111o_1 c261 (.A1(net167),
    .A2(net180),
    .B1(net174),
    .C1(net911),
    .D1(net900),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net171),
    .A1(net183),
    .A2(net181),
    .A3(net112),
    .S0(net911),
    .S1(net806),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net168),
    .A1(net179),
    .A2(net50),
    .A3(net52),
    .S0(net180),
    .S1(net901),
    .X(net185));
 sky130_fd_sc_hd__and2_0 c264 (.A(net74),
    .B(net810),
    .X(net186));
 sky130_fd_sc_hd__and2_1 c265 (.A(net814),
    .B(net64),
    .X(net187));
 sky130_fd_sc_hd__and2_2 c266 (.A(net187),
    .B(net74),
    .X(net188));
 sky130_fd_sc_hd__and2_2 c267 (.A(net186),
    .B(net188),
    .X(net189));
 sky130_fd_sc_hd__and2_2 c268 (.A(net78),
    .B(net188),
    .X(net190));
 sky130_fd_sc_hd__and2_0 c269 (.A(net187),
    .B(net81),
    .X(net191));
 sky130_fd_sc_hd__and3_1 c270 (.A(net188),
    .B(net72),
    .C(net191),
    .X(net192));
 sky130_fd_sc_hd__and2_1 c271 (.A(net188),
    .B(net186),
    .X(net193));
 sky130_fd_sc_hd__and3_1 c272 (.A(net189),
    .B(net79),
    .C(net66),
    .X(net194));
 sky130_fd_sc_hd__and3_2 c273 (.A(net193),
    .B(net188),
    .C(net190),
    .X(net195));
 sky130_fd_sc_hd__and3_2 c274 (.A(net192),
    .B(net194),
    .C(net193),
    .X(net196));
 sky130_fd_sc_hd__and3_1 c275 (.A(net939),
    .B(net191),
    .C(net196),
    .X(net197));
 sky130_fd_sc_hd__and3_1 c276 (.A(net196),
    .B(net189),
    .C(net197),
    .X(net198));
 sky130_fd_sc_hd__and2_1 c277 (.A(net81),
    .B(net196),
    .X(net199));
 sky130_fd_sc_hd__and3_2 c278 (.A(net188),
    .B(net193),
    .C(net933),
    .X(net899));
 sky130_fd_sc_hd__a2111o_2 c279 (.A1(net186),
    .A2(net67),
    .B1(net865),
    .C1(net188),
    .D1(net66),
    .X(net200));
 sky130_fd_sc_hd__and2_1 c280 (.A(net71),
    .B(net76),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net191),
    .A1(net194),
    .A2(net197),
    .A3(net200),
    .S0(net62),
    .S1(net929),
    .X(net202));
 sky130_fd_sc_hd__mux4_2 c282 (.A0(net201),
    .A1(net192),
    .A2(net197),
    .A3(net933),
    .S0(net188),
    .S1(net703),
    .X(net203));
 sky130_fd_sc_hd__and3_1 c283 (.A(net201),
    .B(net200),
    .C(net703),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net187),
    .A1(net204),
    .A2(net939),
    .A3(net190),
    .S0(net197),
    .S1(net860),
    .X(net205));
 sky130_fd_sc_hd__buf_1 c285 (.A(clknet_1_0__leaf_net909),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 c286 (.A(net703),
    .X(net207));
 sky130_fd_sc_hd__and2_1 c287 (.A(net829),
    .B(net807),
    .X(net208));
 sky130_fd_sc_hd__and3_2 c288 (.A(net193),
    .B(net839),
    .C(net208),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c289 (.A(net207),
    .B(net64),
    .C(net839),
    .X(net210));
 sky130_fd_sc_hd__and3_1 c290 (.A(net84),
    .B(net97),
    .C(net192),
    .X(net211));
 sky130_fd_sc_hd__and2_0 c291 (.A(net210),
    .B(net209),
    .X(net212));
 sky130_fd_sc_hd__and3_2 c292 (.A(net74),
    .B(net939),
    .C(net84),
    .X(net213));
 sky130_fd_sc_hd__and2_0 c293 (.A(net212),
    .B(net208),
    .X(net214));
 sky130_fd_sc_hd__and3_1 c294 (.A(net208),
    .B(net213),
    .C(net93),
    .X(net215));
 sky130_fd_sc_hd__and2_0 c295 (.A(net810),
    .B(net204),
    .X(net216));
 sky130_fd_sc_hd__and3_1 c296 (.A(net820),
    .B(net190),
    .C(net213),
    .X(net217));
 sky130_fd_sc_hd__or4bb_1 c297 (.A(net821),
    .B(net211),
    .C_N(net87),
    .D_N(net820),
    .X(net218));
 sky130_fd_sc_hd__and2_1 c298 (.A(net215),
    .B(net860),
    .X(net219));
 sky130_fd_sc_hd__or4bb_1 c299 (.A(net217),
    .B(net216),
    .C_N(net939),
    .D_N(net84),
    .X(net220));
 sky130_fd_sc_hd__a2111o_1 c300 (.A1(net93),
    .A2(net209),
    .B1(net220),
    .C1(net200),
    .D1(net215),
    .X(net221));
 sky130_fd_sc_hd__and3_1 c301 (.A(net219),
    .B(net214),
    .C(net213),
    .X(net222));
 sky130_fd_sc_hd__and2_2 c302 (.A(net210),
    .B(net189),
    .X(net223));
 sky130_fd_sc_hd__or4bb_2 c303 (.A(net220),
    .B(net89),
    .C_N(net223),
    .D_N(net938),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net221),
    .A1(net832),
    .A2(net224),
    .A3(net223),
    .S0(net217),
    .S1(net84),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 c305 (.A(net703),
    .X(net226));
 sky130_fd_sc_hd__sdfrtn_1 c306 (.CLK_N(clknet_4_0_0_clk),
    .D(net218),
    .RESET_B(net219),
    .SCD(net226),
    .SCE(net832),
    .Q(net882));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net214),
    .A1(net225),
    .A2(net990),
    .A3(net226),
    .S0(net209),
    .S1(net223),
    .X(net227));
 sky130_fd_sc_hd__and2_1 c308 (.A(net109),
    .B(net226),
    .X(net228));
 sky130_fd_sc_hd__and2_4 c309 (.A(net117),
    .B(net196),
    .X(net908));
 sky130_fd_sc_hd__buf_1 c310 (.A(net629),
    .X(net229));
 sky130_fd_sc_hd__and2_0 c311 (.A(net824),
    .B(net843),
    .X(net230));
 sky130_fd_sc_hd__and3_1 c312 (.A(net229),
    .B(net3),
    .C(net939),
    .X(net231));
 sky130_fd_sc_hd__and3_2 c313 (.A(net192),
    .B(net189),
    .C(net89),
    .X(net232));
 sky130_fd_sc_hd__or4bb_1 c314 (.A(net205),
    .B(net908),
    .C_N(net209),
    .D_N(net683),
    .X(net233));
 sky130_fd_sc_hd__and3_1 c315 (.A(net231),
    .B(net935),
    .C(net692),
    .X(net234));
 sky130_fd_sc_hd__and2_2 c316 (.A(net64),
    .B(net949),
    .X(net235));
 sky130_fd_sc_hd__or4bb_4 c317 (.A(net87),
    .B(net228),
    .C_N(net89),
    .D_N(net232),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c318 (.A0(net204),
    .A1(net101),
    .A2(net235),
    .A3(net908),
    .S0(net236),
    .S1(net224),
    .X(net237));
 sky130_fd_sc_hd__buf_1 c319 (.A(clknet_1_1__leaf_net909),
    .X(net238));
 sky130_fd_sc_hd__and2_2 c320 (.A(net89),
    .B(net224),
    .X(net239));
 sky130_fd_sc_hd__buf_1 c321 (.A(net629),
    .X(net240));
 sky130_fd_sc_hd__and2_0 c322 (.A(net230),
    .B(net236),
    .X(net241));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net229),
    .A1(net224),
    .A2(net204),
    .A3(net230),
    .S0(net67),
    .S1(net239),
    .X(net242));
 sky130_fd_sc_hd__and3_2 c324 (.A(net231),
    .B(net117),
    .C(net692),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net123),
    .A1(net240),
    .A2(net234),
    .A3(clknet_1_0__leaf_net238),
    .S0(net824),
    .S1(net118),
    .X(net244));
 sky130_fd_sc_hd__and3_1 c326 (.A(clknet_1_1__leaf_net238),
    .B(net115),
    .C(net935),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c327 (.A(net245),
    .B(net882),
    .C(net935),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net241),
    .A1(clknet_1_1__leaf_net246),
    .A2(net235),
    .A3(net224),
    .S0(net935),
    .S1(clknet_1_0__leaf_net718),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net239),
    .A1(clknet_1_0__leaf_net246),
    .A2(net243),
    .A3(net236),
    .S0(net229),
    .S1(clknet_1_1__leaf_net718),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 c330 (.A(net637),
    .X(net249));
 sky130_fd_sc_hd__and2_0 c331 (.A(net249),
    .B(net236),
    .X(net250));
 sky130_fd_sc_hd__and3_1 c332 (.A(net857),
    .B(net226),
    .C(net713),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 c333 (.A(net638),
    .X(net252));
 sky130_fd_sc_hd__and2_2 c334 (.A(net224),
    .B(net127),
    .X(net253));
 sky130_fd_sc_hd__buf_1 c335 (.A(net800),
    .X(net254));
 sky130_fd_sc_hd__and3_1 c336 (.A(net949),
    .B(net254),
    .C(clknet_1_1__leaf_net719),
    .X(net255));
 sky130_fd_sc_hd__buf_1 c337 (.A(net803),
    .X(net892));
 sky130_fd_sc_hd__and3_1 c338 (.A(net209),
    .B(net948),
    .C(net936),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c339 (.A(net939),
    .B(net948),
    .C(net709),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 c340 (.A(net801),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_1 c341 (.A(net712),
    .X(net919));
 sky130_fd_sc_hd__or4bb_1 c342 (.A(net255),
    .B(net929),
    .C_N(net948),
    .D_N(net232),
    .X(net258));
 sky130_fd_sc_hd__and3_1 c343 (.A(net223),
    .B(net938),
    .C(net692),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c344 (.A(net252),
    .B(net134),
    .C(net714),
    .X(net260));
 sky130_fd_sc_hd__or4bb_1 c345 (.A(net232),
    .B(net259),
    .C_N(net254),
    .D_N(net935),
    .X(net261));
 sky130_fd_sc_hd__and2_0 c346 (.A(net259),
    .B(net932),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net796),
    .X(net263));
 sky130_fd_sc_hd__or4bb_1 c348 (.A(net250),
    .B(net932),
    .C_N(net907),
    .D_N(net928),
    .X(net264));
 sky130_fd_sc_hd__a2111o_1 c349 (.A1(net257),
    .A2(net127),
    .B1(net932),
    .C1(net949),
    .D1(clknet_1_0__leaf_net719),
    .X(net265));
 sky130_fd_sc_hd__a2111o_1 c350 (.A1(clknet_1_0__leaf_net265),
    .A2(net932),
    .B1(net928),
    .C1(net679),
    .D1(net692),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net262),
    .A1(clknet_1_1__leaf_net265),
    .A2(net932),
    .A3(net948),
    .S0(net908),
    .S1(net232),
    .X(net267));
 sky130_fd_sc_hd__a2111o_1 c352 (.A1(net256),
    .A2(net914),
    .B1(net936),
    .C1(net908),
    .D1(net709),
    .X(net268));
 sky130_fd_sc_hd__and3_1 c353 (.A(net932),
    .B(net131),
    .C(net716),
    .X(net269));
 sky130_fd_sc_hd__or4bb_4 c354 (.A(net149),
    .B(net835),
    .C_N(net256),
    .D_N(net709),
    .X(net867));
 sky130_fd_sc_hd__sdfbbp_1 c355 (.CLK(clknet_4_4_0_clk),
    .D(net239),
    .RESET_B(net27),
    .SCD(net907),
    .SCE(net154),
    .SET_B(net969),
    .Q(net271),
    .Q_N(net270));
 sky130_fd_sc_hd__and3_1 c356 (.A(net263),
    .B(net867),
    .C(net27),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 c357 (.A(net791),
    .X(net273));
 sky130_fd_sc_hd__and3_1 c358 (.A(net41),
    .B(net939),
    .C(clknet_1_0__leaf_net717),
    .X(net274));
 sky130_fd_sc_hd__and3_1 c359 (.A(net932),
    .B(net682),
    .C(net716),
    .X(net912));
 sky130_fd_sc_hd__or4bb_1 c360 (.A(net27),
    .B(net932),
    .C_N(net263),
    .D_N(net923),
    .X(net275));
 sky130_fd_sc_hd__and3_2 c361 (.A(net932),
    .B(net917),
    .C(net914),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 c362 (.A(net791),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net273),
    .A1(net27),
    .A2(net160),
    .A3(net923),
    .S0(net276),
    .S1(clknet_1_1__leaf_net717),
    .X(net278));
 sky130_fd_sc_hd__buf_2 c364 (.A(net802),
    .X(net885));
 sky130_fd_sc_hd__a2111o_1 c365 (.A1(net885),
    .A2(net149),
    .B1(net898),
    .C1(net867),
    .D1(net725),
    .X(net279));
 sky130_fd_sc_hd__or4bb_2 c366 (.A(net161),
    .B(net882),
    .C_N(net277),
    .D_N(net725),
    .X(net280));
 sky130_fd_sc_hd__buf_1 c367 (.A(net802),
    .X(net281));
 sky130_fd_sc_hd__a2111o_1 c368 (.A1(net277),
    .A2(net281),
    .B1(net885),
    .C1(net261),
    .D1(net724),
    .X(net282));
 sky130_fd_sc_hd__a2111o_1 c369 (.A1(net281),
    .A2(net282),
    .B1(net280),
    .C1(net885),
    .D1(net276),
    .X(net283));
 sky130_fd_sc_hd__sdfbbn_1 c370 (.CLK_N(clknet_4_5_0_clk),
    .D(net280),
    .RESET_B(net279),
    .SCD(net282),
    .SCE(net276),
    .SET_B(clknet_1_1__leaf_net274),
    .Q(net915),
    .Q_N(net284));
 sky130_fd_sc_hd__clkbuf_2 c371 (.A(net799),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net240),
    .A1(net885),
    .A2(net285),
    .A3(net27),
    .S0(net142),
    .S1(net993),
    .X(net286));
 sky130_fd_sc_hd__sdfbbn_2 c373 (.CLK_N(clknet_4_7_0_clk),
    .D(net286),
    .RESET_B(net928),
    .SCD(net912),
    .SCE(net285),
    .SET_B(net976),
    .Q(net893),
    .Q_N(net287));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net279),
    .A1(net181),
    .A2(net911),
    .A3(net923),
    .S0(net912),
    .S1(net893),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net51),
    .A1(net908),
    .A2(net816),
    .A3(net955),
    .S0(net284),
    .S1(net896),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net239),
    .A1(net51),
    .A2(net875),
    .A3(net867),
    .S0(net901),
    .S1(net876),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net818),
    .A1(net174),
    .A2(net907),
    .A3(net912),
    .S0(net896),
    .S1(net876),
    .X(net291));
 sky130_fd_sc_hd__and3_1 c396 (.A(net65),
    .B(net190),
    .C(net939),
    .X(net292));
 sky130_fd_sc_hd__and2_0 c397 (.A(net815),
    .B(clknet_1_0__leaf_net206),
    .X(net293));
 sky130_fd_sc_hd__and2_1 c398 (.A(net67),
    .B(net62),
    .X(net294));
 sky130_fd_sc_hd__or4bb_1 c399 (.A(net811),
    .B(net196),
    .C_N(clknet_1_0__leaf_net293),
    .D_N(net198),
    .X(net295));
 sky130_fd_sc_hd__and2_0 c400 (.A(net294),
    .B(net670),
    .X(net296));
 sky130_fd_sc_hd__sdfbbp_1 c401 (.CLK(clknet_4_0_0_clk),
    .D(net75),
    .RESET_B(net294),
    .SCD(net929),
    .SCE(net194),
    .SET_B(net703),
    .Q(net298),
    .Q_N(net297));
 sky130_fd_sc_hd__or4bb_1 c402 (.A(net813),
    .B(net189),
    .C_N(net194),
    .D_N(net952),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 c403 (.A(net701),
    .X(net300));
 sky130_fd_sc_hd__and2_1 c404 (.A(net807),
    .B(net953),
    .X(net301));
 sky130_fd_sc_hd__and2_0 c405 (.A(clknet_1_0__leaf_net293),
    .B(net296),
    .X(net302));
 sky130_fd_sc_hd__and2_0 c406 (.A(net838),
    .B(net301),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 c407 (.A(net701),
    .X(net304));
 sky130_fd_sc_hd__and2_0 c408 (.A(net197),
    .B(clknet_1_0__leaf_net302),
    .X(net305));
 sky130_fd_sc_hd__sdfbbn_2 c409 (.CLK_N(clknet_4_2_0_clk),
    .D(net294),
    .RESET_B(clknet_1_0__leaf_net305),
    .SCD(net301),
    .SCE(net953),
    .SET_B(net670),
    .Q(net307),
    .Q_N(net306));
 sky130_fd_sc_hd__and3_1 c410 (.A(net292),
    .B(net303),
    .C(net952),
    .X(net308));
 sky130_fd_sc_hd__and2_0 c411 (.A(net308),
    .B(clknet_1_0__leaf_net206),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 c412 (.A(net712),
    .X(net310));
 sky130_fd_sc_hd__or4bb_1 c413 (.A(net301),
    .B(net307),
    .C_N(net310),
    .D_N(net952),
    .X(net311));
 sky130_fd_sc_hd__or4bb_1 c414 (.A(clknet_1_1__leaf_net206),
    .B(net303),
    .C_N(clknet_1_0__leaf_net309),
    .D_N(net952),
    .X(net312));
 sky130_fd_sc_hd__and2_0 c415 (.A(net304),
    .B(net310),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net313),
    .A1(clknet_1_0__leaf_net309),
    .A2(clknet_1_0__leaf_net312),
    .A3(net306),
    .S0(net308),
    .S1(net952),
    .X(net870));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(clknet_1_0__leaf_net305),
    .A1(net313),
    .A2(net307),
    .A3(net308),
    .S0(net310),
    .S1(net952),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 c418 (.A(net665),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net299),
    .A1(net839),
    .A2(clknet_1_0__leaf_net312),
    .A3(net311),
    .S0(net949),
    .S1(net88),
    .X(net316));
 sky130_fd_sc_hd__or4bb_1 c420 (.A(net300),
    .B(net832),
    .C_N(net807),
    .D_N(net223),
    .X(net317));
 sky130_fd_sc_hd__and2_0 c421 (.A(net303),
    .B(net200),
    .X(net318));
 sky130_fd_sc_hd__and2_1 c422 (.A(net865),
    .B(net300),
    .X(net319));
 sky130_fd_sc_hd__and2_1 c423 (.A(net88),
    .B(net319),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 c424 (.A(net665),
    .X(net321));
 sky130_fd_sc_hd__and2_0 c425 (.A(net301),
    .B(clknet_1_1__leaf_net312),
    .X(net322));
 sky130_fd_sc_hd__and3_1 c426 (.A(net321),
    .B(net301),
    .C(net196),
    .X(net323));
 sky130_fd_sc_hd__and2_1 c427 (.A(net96),
    .B(net670),
    .X(net324));
 sky130_fd_sc_hd__and2_0 c428 (.A(net318),
    .B(net323),
    .X(net325));
 sky130_fd_sc_hd__buf_1 c429 (.A(net664),
    .X(net326));
 sky130_fd_sc_hd__and2_1 c430 (.A(net311),
    .B(net310),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net200),
    .A1(net315),
    .A2(net190),
    .A3(net103),
    .S0(net82),
    .S1(net320),
    .X(net328));
 sky130_fd_sc_hd__and3_2 c432 (.A(net317),
    .B(net868),
    .C(net327),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c433 (.A(net92),
    .B(net209),
    .C(net328),
    .X(net330));
 sky130_fd_sc_hd__buf_1 c434 (.A(clknet_1_0__leaf_net794),
    .X(net331));
 sky130_fd_sc_hd__buf_2 c435 (.A(net712),
    .X(net332));
 sky130_fd_sc_hd__and3_1 c436 (.A(net216),
    .B(clknet_1_0__leaf_net331),
    .C(net330),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_4 c437 (.A(net804),
    .X(net890));
 sky130_fd_sc_hd__and3_1 c438 (.A(clknet_1_1__leaf_net331),
    .B(clknet_1_0__leaf_net887),
    .C(net200),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 c439 (.A(net664),
    .X(net334));
 sky130_fd_sc_hd__sdfrtp_4 c440 (.CLK(clknet_4_1_0_clk),
    .D(net243),
    .RESET_B(clknet_1_1__leaf_net887),
    .SCD(net101),
    .SCE(net935),
    .Q(net335));
 sky130_fd_sc_hd__or4bb_1 c441 (.A(net209),
    .B(net115),
    .C_N(net235),
    .D_N(net223),
    .X(net336));
 sky130_fd_sc_hd__or4bb_1 c442 (.A(clknet_1_1__leaf_net293),
    .B(net320),
    .C_N(clknet_1_0__leaf_net333),
    .D_N(net235),
    .X(net337));
 sky130_fd_sc_hd__and3_1 c443 (.A(net805),
    .B(net938),
    .C(net706),
    .X(net338));
 sky130_fd_sc_hd__and3_2 c444 (.A(net953),
    .B(net236),
    .C(net335),
    .X(net879));
 sky130_fd_sc_hd__and3_1 c445 (.A(net338),
    .B(net706),
    .C(net721),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 c446 (.X(net340));
 sky130_fd_sc_hd__buf_1 c447 (.A(net627),
    .X(net341));
 sky130_fd_sc_hd__a2111o_1 c448 (.A1(net82),
    .A2(net336),
    .B1(net929),
    .C1(net341),
    .X(net342));
 sky130_fd_sc_hd__and3_1 c449 (.A(net235),
    .B(net3),
    .C(net320),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net196),
    .A1(net832),
    .A2(net335),
    .A3(net243),
    .S0(net67),
    .S1(net953),
    .X(net344));
 sky130_fd_sc_hd__sdfrtp_4 c451 (.CLK(clknet_4_1_0_clk),
    .D(net118),
    .RESET_B(net235),
    .SCD(net115),
    .SCE(clknet_1_1__leaf_net870),
    .Q(net889));
 sky130_fd_sc_hd__or4bb_4 c452 (.A(net341),
    .B(net889),
    .C_N(net937),
    .D_N(net726),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_1 c453 (.CLK_N(clknet_4_3_0_clk),
    .D(net343),
    .RESET_B(net975),
    .SCD(net934),
    .SCE(clknet_1_0__leaf_net333),
    .SET_B(net981),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__sdfbbp_1 c454 (.CLK(clknet_4_2_0_clk),
    .D(net118),
    .RESET_B(net236),
    .SCD(net934),
    .SCE(net335),
    .SET_B(net726),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net349),
    .A1(net889),
    .A2(net882),
    .A3(clknet_1_0__leaf_net333),
    .S0(net706),
    .S1(net981),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net319),
    .A1(net345),
    .A2(net882),
    .A3(net927),
    .S0(net934),
    .S1(net727),
    .X(net351));
 sky130_fd_sc_hd__mux4_2 c457 (.A0(net115),
    .A1(net223),
    .A2(net346),
    .A3(net934),
    .S0(net335),
    .S1(net727),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net336),
    .A1(net329),
    .A2(net352),
    .A3(net327),
    .S0(net727),
    .S1(net728),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net858),
    .A1(net353),
    .A2(net345),
    .A3(net352),
    .S0(net82),
    .S1(net335),
    .X(net354));
 sky130_fd_sc_hd__sdfbbn_1 c460 (.CLK_N(clknet_4_3_0_clk),
    .D(net338),
    .RESET_B(net353),
    .SCD(net341),
    .SCE(net345),
    .SET_B(net727),
    .Q(net356),
    .Q_N(net355));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net356),
    .A1(net335),
    .A2(net343),
    .A3(net352),
    .S0(net934),
    .S1(net353),
    .X(net357));
 sky130_fd_sc_hd__a2111o_2 c462 (.A1(net327),
    .A2(net377),
    .B1(net372),
    .C1(net335),
    .D1(net733),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net243),
    .A1(net125),
    .A2(net365),
    .A3(net670),
    .S0(net731),
    .S1(net733),
    .X(net359));
 sky130_fd_sc_hd__or4bb_1 c464 (.A(net369),
    .B(net373),
    .C_N(net378),
    .D_N(net358),
    .X(net360));
 sky130_fd_sc_hd__a2111o_1 c465 (.A1(net189),
    .A2(net889),
    .B1(clknet_1_0__leaf_net360),
    .C1(net365),
    .D1(net968),
    .X(net361));
 sky130_fd_sc_hd__sdfbbn_1 c466 (.CLK_N(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net360),
    .RESET_B(clknet_1_1__leaf_net333),
    .SCD(net371),
    .SCE(net874),
    .SET_B(net667),
    .Q(net363),
    .Q_N(net362));
 sky130_fd_sc_hd__a2111o_1 c467 (.A1(net345),
    .A2(net372),
    .B1(net378),
    .C1(net667),
    .D1(net733),
    .X(net902));
 sky130_fd_sc_hd__and3_1 c468 (.A(net136),
    .B(net949),
    .C(net723),
    .X(net364));
 sky130_fd_sc_hd__buf_2 c469 (.A(net988),
    .X(net365));
 sky130_fd_sc_hd__and3_1 c470 (.A(net332),
    .B(net335),
    .C(net868),
    .X(net366));
 sky130_fd_sc_hd__and3_1 c471 (.A(net366),
    .B(net3),
    .C(net948),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 c472 (.A(net988),
    .X(net368));
 sky130_fd_sc_hd__buf_1 c473 (.A(clknet_1_1__leaf_net793),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 c474 (.A(net801),
    .X(net370));
 sky130_fd_sc_hd__or4bb_2 c475 (.A(net236),
    .B(net223),
    .C_N(net92),
    .D_N(net729),
    .X(net371));
 sky130_fd_sc_hd__or4bb_2 c476 (.A(net368),
    .B(net370),
    .C_N(net937),
    .D_N(net730),
    .X(net372));
 sky130_fd_sc_hd__sdfrtp_2 c477 (.CLK(clknet_4_3_0_clk),
    .D(net370),
    .RESET_B(net236),
    .SCD(net927),
    .SCE(net366),
    .Q(net373));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net125),
    .A1(net372),
    .A2(net134),
    .A3(net373),
    .S0(net243),
    .S1(net335),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net372),
    .A1(net243),
    .A2(clknet_1_0__leaf_net333),
    .A3(net710),
    .S0(net730),
    .S1(net732),
    .X(net375));
 sky130_fd_sc_hd__buf_1 c480 (.A(net803),
    .X(net886));
 sky130_fd_sc_hd__a2111o_4 c481 (.A1(net223),
    .A2(net948),
    .B1(net143),
    .C1(net723),
    .D1(net732),
    .X(net874));
 sky130_fd_sc_hd__sdfbbp_1 c482 (.CLK(clknet_4_6_0_clk),
    .D(net368),
    .RESET_B(net874),
    .SCD(clknet_1_1__leaf_net333),
    .SCE(net987),
    .SET_B(net968),
    .Q(net377),
    .Q_N(net376));
 sky130_fd_sc_hd__a2111o_2 c483 (.A1(net838),
    .A2(net372),
    .B1(net373),
    .C1(net949),
    .D1(net734),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net165),
    .A1(net276),
    .A2(net948),
    .A3(net41),
    .S0(net287),
    .S1(net895),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net276),
    .A1(net165),
    .A2(net948),
    .A3(net937),
    .S0(net927),
    .S1(net42),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net143),
    .A1(net885),
    .A2(net271),
    .A3(net948),
    .S0(net35),
    .S1(clknet_1_0__leaf_net736),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net269),
    .A1(net376),
    .A2(clknet_1_0__leaf_net381),
    .A3(net287),
    .S0(net895),
    .S1(net884),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net358),
    .A1(net874),
    .A2(net893),
    .A3(net149),
    .S0(net885),
    .S1(net270),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net383),
    .A1(clknet_1_0__leaf_net381),
    .A2(net346),
    .A3(net269),
    .S0(clknet_1_1__leaf_net887),
    .S1(net358),
    .X(net384));
 sky130_fd_sc_hd__mux4_2 c490 (.A0(net36),
    .A1(net270),
    .A2(net41),
    .A3(net376),
    .S0(net666),
    .S1(clknet_1_1__leaf_net736),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(clknet_1_0__leaf_net925),
    .A1(net285),
    .A2(net358),
    .A3(clknet_1_1__leaf_net333),
    .S0(net893),
    .S1(net666),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net41),
    .A1(net165),
    .A2(clknet_1_1__leaf_net333),
    .A3(net383),
    .S0(clknet_1_0__leaf_net736),
    .S1(clknet_1_0__leaf_net737),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net347),
    .A1(net276),
    .A2(net927),
    .A3(net735),
    .S0(clknet_1_0__leaf_net897),
    .S1(net741),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(clknet_1_1__leaf_net333),
    .A1(net902),
    .A2(net885),
    .A3(net715),
    .S0(clknet_1_0__leaf_net737),
    .S1(net740),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net269),
    .A1(net285),
    .A2(net895),
    .A3(clknet_1_0__leaf_net897),
    .S0(clknet_1_1__leaf_net737),
    .S1(net740),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net335),
    .A1(net886),
    .A2(net929),
    .A3(net165),
    .S0(net738),
    .S1(net891),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net371),
    .A1(net165),
    .A2(net735),
    .A3(clknet_1_1__leaf_net736),
    .S0(net741),
    .S1(net742),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net890),
    .A1(net35),
    .A2(net287),
    .A3(net735),
    .S0(net742),
    .S1(net744),
    .X(net392));
 sky130_fd_sc_hd__sdfbbn_1 c499 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net925),
    .RESET_B(clknet_1_1__leaf_net333),
    .SCD(clknet_1_1__leaf_net381),
    .SCE(net903),
    .SET_B(net744),
    .Q(net394),
    .Q_N(net393));
 sky130_fd_sc_hd__mux4_2 c500 (.A0(net285),
    .A1(net36),
    .A2(net938),
    .A3(net738),
    .S0(net743),
    .S1(net744),
    .X(net395));
 sky130_fd_sc_hd__mux4_2 c501 (.A0(net392),
    .A1(net880),
    .A2(net395),
    .A3(net285),
    .S0(net891),
    .S1(net744),
    .X(net866));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net276),
    .A1(net395),
    .A2(net393),
    .A3(net971),
    .S0(net995),
    .S1(net744),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 c503 (.A0(net35),
    .A1(clknet_1_1__leaf_net381),
    .A2(clknet_1_0__leaf_net925),
    .A3(net395),
    .S0(net738),
    .S1(net744),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net347),
    .A1(net394),
    .A2(net253),
    .A3(clknet_1_1__leaf_net397),
    .S0(net937),
    .S1(net744),
    .X(net398));
 sky130_fd_sc_hd__mux4_2 c505 (.A0(net134),
    .A1(clknet_1_0__leaf_net397),
    .A2(net285),
    .A3(net892),
    .S0(net395),
    .S1(net744),
    .X(net399));
 sky130_fd_sc_hd__and3_1 c528 (.A(net200),
    .B(net190),
    .C(net75),
    .X(net400));
 sky130_fd_sc_hd__and2_2 c529 (.A(net815),
    .B(net66),
    .X(net401));
 sky130_fd_sc_hd__and3_2 c530 (.A(net308),
    .B(net401),
    .C(net952),
    .X(net402));
 sky130_fd_sc_hd__and3_2 c531 (.A(net813),
    .B(net307),
    .C(net310),
    .X(net403));
 sky130_fd_sc_hd__buf_2 c532 (.A(net688),
    .X(net404));
 sky130_fd_sc_hd__and3_1 c533 (.A(net307),
    .B(net400),
    .C(net402),
    .X(net405));
 sky130_fd_sc_hd__and3_1 c534 (.A(net405),
    .B(net404),
    .C(net66),
    .X(net406));
 sky130_fd_sc_hd__and2_1 c535 (.A(net194),
    .B(net405),
    .X(net407));
 sky130_fd_sc_hd__buf_1 c536 (.A(net688),
    .X(net408));
 sky130_fd_sc_hd__buf_1 c537 (.A(net653),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 c538 (.A(net687),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 c539 (.A(net650),
    .X(net411));
 sky130_fd_sc_hd__sdfsbp_1 c540 (.CLK(clknet_4_8_0_clk),
    .D(net407),
    .SCD(net813),
    .SCE(net410),
    .SET_B(net944),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__mux4_2 c541 (.A0(net62),
    .A1(net413),
    .A2(net409),
    .A3(net402),
    .S0(net306),
    .S1(net944),
    .X(net414));
 sky130_fd_sc_hd__a2111o_1 c542 (.A1(net400),
    .A2(net307),
    .B1(net409),
    .C1(net412),
    .D1(net944),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 c543 (.A0(net415),
    .A1(net408),
    .A2(net401),
    .A3(net400),
    .S0(net306),
    .S1(net953),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net404),
    .A1(net414),
    .A2(net412),
    .A3(net944),
    .S0(net410),
    .S1(net952),
    .X(net417));
 sky130_fd_sc_hd__sdfbbn_1 c545 (.CLK_N(clknet_4_8_0_clk),
    .D(net409),
    .RESET_B(net416),
    .SCD(net417),
    .SCE(net944),
    .SET_B(net297),
    .Q(net419),
    .Q_N(net418));
 sky130_fd_sc_hd__mux4_1 c546 (.A0(net417),
    .A1(net419),
    .A2(net415),
    .A3(net403),
    .S0(net412),
    .S1(net944),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net419),
    .A1(net414),
    .A2(net415),
    .A3(net308),
    .S0(net417),
    .S1(net745),
    .X(net421));
 sky130_fd_sc_hd__mux4_2 c548 (.A0(net413),
    .A1(net944),
    .A2(net418),
    .A3(net402),
    .S0(net745),
    .S1(net746),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net408),
    .A1(net422),
    .A2(net401),
    .A3(net414),
    .S0(net745),
    .S1(net746),
    .X(net423));
 sky130_fd_sc_hd__and3_1 c550 (.A(net326),
    .B(net400),
    .C(net328),
    .X(net424));
 sky130_fd_sc_hd__buf_1 c551 (.A(net702),
    .X(net425));
 sky130_fd_sc_hd__and3_1 c552 (.A(net324),
    .B(net422),
    .C(net945),
    .X(net426));
 sky130_fd_sc_hd__mux4_2 c553 (.A0(net190),
    .A1(net310),
    .A2(net414),
    .A3(net890),
    .S0(net422),
    .S1(net945),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net414),
    .A1(net329),
    .A2(net334),
    .A3(net816),
    .S0(net933),
    .S1(net416),
    .X(net428));
 sky130_fd_sc_hd__sdfsbp_1 c555 (.CLK(clknet_4_8_0_clk),
    .D(net428),
    .SCD(net103),
    .SCE(net427),
    .SET_B(net933),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__or4bb_4 c556 (.A(net328),
    .B(net403),
    .C_N(net401),
    .D_N(net226),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c557 (.A(net330),
    .B(net402),
    .C(net424),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net323),
    .A1(net310),
    .A2(net429),
    .A3(net425),
    .S0(net326),
    .S1(net945),
    .X(net433));
 sky130_fd_sc_hd__buf_1 c559 (.A(net702),
    .X(net434));
 sky130_fd_sc_hd__sdfstp_2 c560 (.CLK(clknet_4_9_0_clk),
    .D(net222),
    .SCD(net992),
    .SCE(net427),
    .SET_B(net974),
    .Q(net435));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(net325),
    .A1(net433),
    .A2(net431),
    .A3(net943),
    .S0(net944),
    .S1(net297),
    .X(net436));
 sky130_fd_sc_hd__and3_1 c562 (.A(net424),
    .B(net943),
    .C(net747),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net432),
    .A1(net943),
    .A2(net832),
    .A3(net403),
    .S0(net404),
    .S1(net435),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net427),
    .A1(net401),
    .A2(net402),
    .A3(net435),
    .S0(net416),
    .S1(net945),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net438),
    .A1(net435),
    .A2(net437),
    .A3(net422),
    .S0(net943),
    .S1(net747),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net628),
    .A1(net222),
    .A2(net432),
    .A3(net435),
    .S0(net427),
    .S1(net747),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c567 (.A(net945),
    .B(net668),
    .C(net747),
    .X(net442));
 sky130_fd_sc_hd__and3_4 c568 (.A(net442),
    .B(net330),
    .C(net422),
    .X(net872));
 sky130_fd_sc_hd__sdfstp_1 c569 (.CLK(clknet_4_8_0_clk),
    .D(net433),
    .SCD(net428),
    .SCE(clknet_1_0__leaf_net870),
    .SET_B(net973),
    .Q(net443));
 sky130_fd_sc_hd__sdfstp_1 c570 (.CLK(clknet_4_9_0_clk),
    .D(net438),
    .SCD(net404),
    .SCE(net435),
    .SET_B(net967),
    .Q(net444));
 sky130_fd_sc_hd__sdfbbp_1 c571 (.CLK(clknet_4_9_0_clk),
    .D(net400),
    .RESET_B(net872),
    .SCD(net994),
    .SCE(net431),
    .SET_B(net945),
    .Q(net446),
    .Q_N(net445));
 sky130_fd_sc_hd__a2111o_1 c572 (.A1(net446),
    .A2(net352),
    .B1(net839),
    .C1(net728),
    .D1(net747),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 c573 (.A(net693),
    .X(net448));
 sky130_fd_sc_hd__sedfxbp_1 c574 (.CLK(clknet_4_9_0_clk),
    .D(net447),
    .DE(net329),
    .SCD(net943),
    .SCE(net835),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__and3_2 c575 (.A(net437),
    .B(net450),
    .C(net745),
    .X(net451));
 sky130_fd_sc_hd__a2111o_1 c576 (.A1(net448),
    .A2(net101),
    .B1(net416),
    .C1(net329),
    .D1(net431),
    .X(net452));
 sky130_fd_sc_hd__or4bb_4 c577 (.A(net450),
    .B(net937),
    .C_N(net352),
    .D_N(net947),
    .X(net453));
 sky130_fd_sc_hd__and3_1 c578 (.A(net832),
    .B(net356),
    .C(net745),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net693),
    .X(net455));
 sky130_fd_sc_hd__and3_2 c580 (.A(net431),
    .B(net832),
    .C(net721),
    .X(net456));
 sky130_fd_sc_hd__and3_1 c581 (.A(net454),
    .B(net450),
    .C(net456),
    .X(net457));
 sky130_fd_sc_hd__and3_1 c582 (.A(net443),
    .B(net451),
    .C(net456),
    .X(net458));
 sky130_fd_sc_hd__a2111o_1 c583 (.A1(net425),
    .A2(net839),
    .B1(net453),
    .C1(net451),
    .D1(net979),
    .X(net459));
 sky130_fd_sc_hd__and3_1 c584 (.A(net456),
    .B(net673),
    .C(net720),
    .X(net460));
 sky130_fd_sc_hd__and3_2 c585 (.A(net320),
    .B(net460),
    .C(net443),
    .X(net461));
 sky130_fd_sc_hd__buf_1 c586 (.A(clknet_1_0__leaf_net793),
    .X(net462));
 sky130_fd_sc_hd__and3_1 c587 (.A(net462),
    .B(net868),
    .C(net931),
    .X(net463));
 sky130_fd_sc_hd__sdfbbn_1 c588 (.CLK_N(clknet_4_9_0_clk),
    .D(net425),
    .RESET_B(net461),
    .SCD(net456),
    .SCE(clknet_1_0__leaf_net870),
    .SET_B(net980),
    .Q(net465),
    .Q_N(net464));
 sky130_fd_sc_hd__sdfbbn_1 c589 (.CLK_N(clknet_4_9_0_clk),
    .D(net982),
    .RESET_B(net890),
    .SCD(net453),
    .SCE(net931),
    .SET_B(net980),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__a2111o_1 c590 (.A1(net226),
    .A2(net466),
    .B1(net454),
    .C1(net817),
    .D1(net728),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net329),
    .A1(net467),
    .A2(net832),
    .A3(net451),
    .S0(net453),
    .S1(net693),
    .X(net469));
 sky130_fd_sc_hd__mux4_2 c592 (.A0(net352),
    .A1(net451),
    .A2(net437),
    .A3(net456),
    .S0(net673),
    .S1(net731),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net468),
    .A1(net467),
    .A2(net470),
    .A3(net449),
    .S0(net464),
    .S1(net748),
    .X(net471));
 sky130_fd_sc_hd__sdfbbp_1 c594 (.CLK(clknet_4_12_0_clk),
    .D(net984),
    .RESET_B(net928),
    .SCD(net872),
    .SCE(net960),
    .SET_B(net977),
    .Q(net473),
    .Q_N(net472));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(clknet_1_1__leaf_net870),
    .A1(net860),
    .A2(net872),
    .A3(net843),
    .S0(net431),
    .S1(net710),
    .X(net474));
 sky130_fd_sc_hd__a2111o_1 c596 (.A1(net435),
    .A2(net960),
    .B1(net378),
    .C1(net416),
    .D1(net937),
    .X(net475));
 sky130_fd_sc_hd__or4bb_1 c597 (.A(net808),
    .B(net931),
    .C_N(net937),
    .D_N(net748),
    .X(net476));
 sky130_fd_sc_hd__a2111o_1 c598 (.A1(net363),
    .A2(net404),
    .B1(net226),
    .C1(net947),
    .D1(net668),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net226),
    .A1(net199),
    .A2(net872),
    .A3(net416),
    .S0(net949),
    .S1(net947),
    .X(net478));
 sky130_fd_sc_hd__sdfbbn_1 c600 (.CLK_N(clknet_4_3_0_clk),
    .D(net404),
    .RESET_B(net365),
    .SCD(net860),
    .SCE(net928),
    .SET_B(net749),
    .Q(net480),
    .Q_N(net479));
 sky130_fd_sc_hd__sdfbbn_1 c601 (.CLK_N(clknet_4_12_0_clk),
    .D(net455),
    .RESET_B(net978),
    .SCD(net101),
    .SCE(net373),
    .SET_B(net416),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net431),
    .A1(net479),
    .A2(net872),
    .A3(net466),
    .S0(net376),
    .S1(net749),
    .X(net483));
 sky130_fd_sc_hd__a2111o_2 c603 (.A1(net960),
    .A2(net482),
    .B1(net839),
    .C1(net435),
    .D1(net835),
    .X(net926));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net373),
    .A1(net482),
    .A2(net928),
    .A3(net456),
    .S0(net874),
    .S1(net693),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net860),
    .A1(net358),
    .A2(net435),
    .A3(net362),
    .S0(net475),
    .S1(net991),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net431),
    .A1(net17),
    .A2(net874),
    .A3(net479),
    .S0(net668),
    .S1(net676),
    .X(net486));
 sky130_fd_sc_hd__a2111o_1 c607 (.A1(net816),
    .A2(net942),
    .B1(net835),
    .C1(net732),
    .D1(net753),
    .X(net487));
 sky130_fd_sc_hd__sdfbbp_1 c608 (.CLK(clknet_4_6_0_clk),
    .D(net486),
    .RESET_B(net927),
    .SCD(net226),
    .SCE(net933),
    .SET_B(net942),
    .Q(net489),
    .Q_N(net488));
 sky130_fd_sc_hd__mux4_2 c609 (.A0(net817),
    .A1(net843),
    .A2(net942),
    .A3(net455),
    .S0(net752),
    .S1(net753),
    .X(net873));
 sky130_fd_sc_hd__a2111o_4 c610 (.A1(net416),
    .A2(net873),
    .B1(net486),
    .C1(net942),
    .D1(net937),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net345),
    .A1(net934),
    .A2(net487),
    .A3(net481),
    .S0(net490),
    .S1(net942),
    .X(net491));
 sky130_fd_sc_hd__a2111o_1 c612 (.A1(net491),
    .A2(net490),
    .B1(net873),
    .C1(net942),
    .D1(net752),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net475),
    .A1(net492),
    .A2(net480),
    .A3(net491),
    .S0(net481),
    .S1(net226),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net487),
    .A1(net477),
    .A2(net873),
    .A3(net491),
    .S0(net942),
    .S1(net748),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net494),
    .A1(net472),
    .A2(net491),
    .A3(net704),
    .S0(net749),
    .S1(net985),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net149),
    .A1(net489),
    .A2(net942),
    .A3(net939),
    .S0(net874),
    .S1(net872),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net377),
    .A1(net867),
    .A2(net927),
    .A3(clknet_1_1__leaf_net925),
    .S0(net921),
    .S1(net866),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net271),
    .A1(net377),
    .A2(net867),
    .A3(clknet_1_0__leaf_net399),
    .S0(net253),
    .S1(net843),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net363),
    .A1(net930),
    .A2(net928),
    .A3(net927),
    .S0(clknet_1_1__leaf_net399),
    .S1(clknet_1_0__leaf_net755),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c62 (.A0(net862),
    .A1(net843),
    .A2(net853),
    .A3(net845),
    .S0(net852),
    .S1(net856),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net928),
    .A1(net358),
    .A2(net927),
    .A3(clknet_1_0__leaf_net399),
    .S0(net942),
    .S1(net131),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net933),
    .A1(net451),
    .A2(net942),
    .A3(clknet_1_0__leaf_net399),
    .S0(net939),
    .S1(clknet_1_0__leaf_net757),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net195),
    .A1(net395),
    .A2(net927),
    .A3(net890),
    .S0(net867),
    .S1(net739),
    .X(net502));
 sky130_fd_sc_hd__mux4_2 c623 (.A0(net42),
    .A1(net451),
    .A2(net149),
    .A3(net395),
    .S0(net488),
    .S1(net378),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net873),
    .A1(net890),
    .A2(net503),
    .A3(net879),
    .S0(net866),
    .S1(net700),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net131),
    .A1(net921),
    .A2(net937),
    .A3(net873),
    .S0(net872),
    .S1(net739),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net503),
    .A1(net36),
    .A2(net872),
    .A3(net868),
    .S0(net695),
    .S1(clknet_1_0__leaf_net757),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net36),
    .A1(net921),
    .A2(net503),
    .A3(net938),
    .S0(net739),
    .S1(clknet_1_0__leaf_net756),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net921),
    .A1(net488),
    .A2(clknet_1_1__leaf_net870),
    .A3(net677),
    .S0(net762),
    .S1(net877),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net378),
    .A1(clknet_1_1__leaf_net870),
    .A2(net930),
    .A3(net761),
    .S0(net877),
    .S1(net763),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net840),
    .A1(net865),
    .A2(net859),
    .A3(net855),
    .S0(net845),
    .S1(net843),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net874),
    .A1(net926),
    .A2(net875),
    .A3(net705),
    .S0(net762),
    .S1(net877),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net451),
    .A1(clknet_1_1__leaf_net870),
    .A2(net956),
    .A3(net708),
    .S0(net739),
    .S1(net763),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_1__leaf_net399),
    .A1(net931),
    .A2(net510),
    .A3(net451),
    .S0(net131),
    .S1(net711),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net878),
    .A1(net867),
    .A2(clknet_1_1__leaf_net757),
    .A3(net761),
    .S0(net763),
    .S1(net764),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net131),
    .A1(net503),
    .A2(net707),
    .A3(net758),
    .S0(net760),
    .S1(net986),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net510),
    .A1(net378),
    .A2(net921),
    .A3(clknet_1_1__leaf_net399),
    .S0(net763),
    .S1(net765),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net513),
    .A1(net377),
    .A2(net866),
    .A3(net677),
    .S0(net877),
    .S1(net764),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net843),
    .A1(net510),
    .A2(clknet_1_1__leaf_net757),
    .A3(net764),
    .S0(net766),
    .S1(net767),
    .X(net517));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net845),
    .A1(net852),
    .A2(net840),
    .A3(net0),
    .S0(net856),
    .S1(net857),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net848),
    .A1(net836),
    .A2(net830),
    .A3(net850),
    .S0(net856),
    .S1(net847),
    .X(net3));
 sky130_fd_sc_hd__a2111o_1 c66 (.A1(net838),
    .A2(net831),
    .B1(net16),
    .C1(net918),
    .D1(net20),
    .X(net4));
 sky130_fd_sc_hd__and2_0 c660 (.A(net80),
    .B(net808),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 c661 (.A(net685),
    .X(net519));
 sky130_fd_sc_hd__buf_1 c662 (.A(net685),
    .X(net520));
 sky130_fd_sc_hd__buf_1 c663 (.A(net652),
    .X(net521));
 sky130_fd_sc_hd__and2_2 c664 (.A(net66),
    .B(net953),
    .X(net522));
 sky130_fd_sc_hd__or4bb_1 c665 (.A(net188),
    .B(net423),
    .C_N(net406),
    .D_N(net412),
    .X(net523));
 sky130_fd_sc_hd__and2_0 c666 (.A(net953),
    .B(net521),
    .X(net524));
 sky130_fd_sc_hd__and2_2 c667 (.A(net402),
    .B(net519),
    .X(net525));
 sky130_fd_sc_hd__or4bb_2 c668 (.A(net413),
    .B(net518),
    .C_N(net525),
    .D_N(net521),
    .X(net526));
 sky130_fd_sc_hd__and2_1 c669 (.A(net518),
    .B(net746),
    .X(net527));
 sky130_fd_sc_hd__and2_0 c67 (.A(net21),
    .B(net20),
    .X(net5));
 sky130_fd_sc_hd__and2_0 c670 (.A(net75),
    .B(net525),
    .X(net528));
 sky130_fd_sc_hd__buf_1 c671 (.A(net651),
    .X(net529));
 sky130_fd_sc_hd__and2_0 c672 (.A(net527),
    .B(net686),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_2 c673 (.A(net687),
    .X(net531));
 sky130_fd_sc_hd__and2_0 c674 (.A(net408),
    .B(net953),
    .X(net532));
 sky130_fd_sc_hd__and3_2 c675 (.A(net72),
    .B(net520),
    .C(net527),
    .X(net533));
 sky130_fd_sc_hd__and3_1 c676 (.A(net410),
    .B(net525),
    .C(net953),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(net532),
    .A1(net522),
    .A2(net531),
    .A3(net406),
    .S0(net534),
    .S1(net80),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net530),
    .A1(net531),
    .A2(net527),
    .A3(net66),
    .S0(net413),
    .S1(net188),
    .X(net536));
 sky130_fd_sc_hd__and3_1 c679 (.A(net536),
    .B(net808),
    .C(net769),
    .X(net537));
 sky130_fd_sc_hd__and2_4 c68 (.A(net20),
    .B(net814),
    .X(net6));
 sky130_fd_sc_hd__and3_1 c680 (.A(net532),
    .B(net946),
    .C(net769),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net521),
    .A1(net538),
    .A2(net533),
    .A3(net536),
    .S0(net686),
    .S1(net768),
    .X(net539));
 sky130_fd_sc_hd__buf_1 c682 (.A(clknet_1_0__leaf_net792),
    .X(net540));
 sky130_fd_sc_hd__and3_1 c683 (.A(clknet_1_0__leaf_net540),
    .B(net818),
    .C(net539),
    .X(net541));
 sky130_fd_sc_hd__and3_1 c684 (.A(net524),
    .B(net444),
    .C(net953),
    .X(net542));
 sky130_fd_sc_hd__and3_1 c685 (.A(net401),
    .B(net298),
    .C(net70),
    .X(net543));
 sky130_fd_sc_hd__and3_1 c686 (.A(net403),
    .B(clknet_1_1__leaf_net540),
    .C(net434),
    .X(net544));
 sky130_fd_sc_hd__buf_1 c687 (.A(clknet_1_1__leaf_net792),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 c688 (.A(net712),
    .X(net546));
 sky130_fd_sc_hd__and3_1 c689 (.A(net430),
    .B(net422),
    .C(net401),
    .X(net547));
 sky130_fd_sc_hd__and3_4 c69 (.A(net6),
    .B(net15),
    .C(net16),
    .X(net7));
 sky130_fd_sc_hd__buf_2 c690 (.A(net798),
    .X(net548));
 sky130_fd_sc_hd__and3_2 c691 (.A(net538),
    .B(net546),
    .C(net531),
    .X(net549));
 sky130_fd_sc_hd__buf_1 c692 (.A(net804),
    .X(net550));
 sky130_fd_sc_hd__buf_1 c693 (.A(net797),
    .X(net551));
 sky130_fd_sc_hd__sdfbbn_1 c694 (.CLK_N(clknet_4_10_0_clk),
    .D(net547),
    .RESET_B(net546),
    .SCD(net537),
    .SCE(net941),
    .SET_B(net543),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__or4bb_1 c695 (.A(net528),
    .B(net941),
    .C_N(net534),
    .D_N(net542),
    .X(net554));
 sky130_fd_sc_hd__a2111o_1 c696 (.A1(net545),
    .A2(net553),
    .B1(net526),
    .C1(net941),
    .D1(net522),
    .X(net555));
 sky130_fd_sc_hd__a2111o_1 c697 (.A1(net544),
    .A2(net941),
    .B1(net552),
    .C1(net527),
    .D1(net691),
    .X(net556));
 sky130_fd_sc_hd__and3_2 c698 (.A(net543),
    .B(net941),
    .C(net553),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net213),
    .A1(net557),
    .A2(net552),
    .A3(net941),
    .S0(net547),
    .S1(net691),
    .X(net558));
 sky130_fd_sc_hd__and3_4 c70 (.A(net7),
    .B(net6),
    .C(net4),
    .X(net880));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net527),
    .A1(net553),
    .A2(net557),
    .A3(net941),
    .S0(net546),
    .S1(net770),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net559),
    .A1(net553),
    .A2(clknet_1_0__leaf_net556),
    .A3(net557),
    .S0(net298),
    .S1(net941),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net560),
    .A1(net539),
    .A2(net524),
    .A3(net941),
    .S0(net552),
    .S1(net770),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net444),
    .A1(clknet_1_0__leaf_net556),
    .A2(net401),
    .A3(clknet_1_0__leaf_net561),
    .S0(net332),
    .S1(net557),
    .X(net562));
 sky130_fd_sc_hd__a2111o_1 c704 (.A1(net538),
    .A2(net103),
    .B1(net461),
    .C1(net298),
    .D1(net770),
    .X(net563));
 sky130_fd_sc_hd__a2111o_1 c705 (.A1(net550),
    .A2(net461),
    .B1(clknet_1_0__leaf_net556),
    .C1(net538),
    .D1(net938),
    .X(net564));
 sky130_fd_sc_hd__a2111o_4 c706 (.A1(net529),
    .A2(net557),
    .B1(net550),
    .C1(net931),
    .D1(net770),
    .X(net565));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_11_0_clk),
    .D(net563),
    .RESET_B(net461),
    .SCD(net549),
    .SCE(net933),
    .SET_B(net989),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__buf_1 c708 (.A(clknet_1_1__leaf_net794),
    .X(net568));
 sky130_fd_sc_hd__or4bb_1 c709 (.A(net520),
    .B(net565),
    .C_N(clknet_1_0__leaf_net568),
    .D_N(net931),
    .X(net569));
 sky130_fd_sc_hd__or4bb_1 c71 (.A(net6),
    .B(net862),
    .C_N(net950),
    .D_N(net880),
    .X(net8));
 sky130_fd_sc_hd__a2111o_1 c710 (.A1(net946),
    .A2(net520),
    .B1(clknet_1_0__leaf_net556),
    .C1(net690),
    .D1(net771),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(clknet_1_1__leaf_net561),
    .A1(net546),
    .A2(net565),
    .A3(net461),
    .S0(net946),
    .S1(net943),
    .X(net571));
 sky130_fd_sc_hd__sdfbbp_1 c712 (.CLK(clknet_4_14_0_clk),
    .D(net463),
    .RESET_B(net565),
    .SCD(net456),
    .SCE(net101),
    .SET_B(net970),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__sdfbbn_2 c713 (.CLK_N(clknet_4_11_0_clk),
    .D(net998),
    .RESET_B(net817),
    .SCD(net943),
    .SCE(net565),
    .SET_B(net102),
    .Q(net575),
    .Q_N(net574));
 sky130_fd_sc_hd__a2111o_1 c714 (.A1(net531),
    .A2(net808),
    .B1(net565),
    .C1(net533),
    .D1(net411),
    .X(net576));
 sky130_fd_sc_hd__a2111o_1 c715 (.A1(net457),
    .A2(clknet_1_0__leaf_net556),
    .B1(net298),
    .C1(net461),
    .D1(net931),
    .X(net577));
 sky130_fd_sc_hd__a2111o_4 c716 (.A1(net557),
    .A2(net548),
    .B1(net566),
    .C1(net574),
    .D1(net751),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net564),
    .A1(net103),
    .A2(net933),
    .A3(net525),
    .S0(net101),
    .S1(clknet_1_0__leaf_net699),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net570),
    .A1(net577),
    .A2(net332),
    .A3(net578),
    .S0(net944),
    .S1(net349),
    .X(net580));
 sky130_fd_sc_hd__a2111o_2 c719 (.A1(net573),
    .A2(net578),
    .B1(net934),
    .C1(net678),
    .D1(net770),
    .X(net581));
 sky130_fd_sc_hd__a2111o_4 c72 (.A1(net7),
    .A2(net950),
    .B1(net16),
    .C1(net23),
    .D1(net850),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_1__leaf_net568),
    .A1(net943),
    .A2(net581),
    .A3(net565),
    .S0(net548),
    .S1(clknet_1_0__leaf_net773),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net529),
    .A1(net581),
    .A2(net578),
    .A3(net678),
    .S0(net772),
    .S1(clknet_1_1__leaf_net773),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net943),
    .A1(net572),
    .A2(clknet_1_1__leaf_net583),
    .A3(net578),
    .S0(net751),
    .S1(clknet_1_0__leaf_net774),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net537),
    .A1(clknet_1_0__leaf_net583),
    .A2(net946),
    .A3(net581),
    .S0(net771),
    .S1(clknet_1_0__leaf_net775),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_0__leaf_net583),
    .A1(net578),
    .A2(net581),
    .A3(net934),
    .S0(clknet_1_0__leaf_net775),
    .S1(net777),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net567),
    .A1(net581),
    .A2(net549),
    .A3(clknet_1_1__leaf_net775),
    .S0(net776),
    .S1(net778),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net101),
    .A1(net522),
    .A2(net578),
    .A3(net947),
    .S0(net938),
    .S1(net70),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net467),
    .A1(net565),
    .A2(net473),
    .A3(net332),
    .S0(net546),
    .S1(clknet_1_0__leaf_net755),
    .X(net589));
 sky130_fd_sc_hd__a2111o_1 c728 (.A1(net816),
    .A2(net533),
    .B1(net772),
    .C1(clknet_1_1__leaf_net774),
    .D1(net780),
    .X(net590));
 sky130_fd_sc_hd__a2111o_1 c729 (.A1(net456),
    .A2(net817),
    .B1(net549),
    .C1(net578),
    .D1(clknet_1_0__leaf_net774),
    .X(net591));
 sky130_fd_sc_hd__and2_0 c73 (.A(net9),
    .B(net821),
    .X(net10));
 sky130_fd_sc_hd__a2111o_1 c730 (.A1(net581),
    .A2(net549),
    .B1(net533),
    .C1(net578),
    .D1(net476),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net470),
    .A1(net934),
    .A2(net581),
    .A3(clknet_1_0__leaf_net591),
    .S0(net574),
    .S1(net779),
    .X(net593));
 sky130_fd_sc_hd__sdfbbn_2 c732 (.CLK_N(clknet_4_14_0_clk),
    .D(net476),
    .RESET_B(net565),
    .SCD(clknet_1_0__leaf_net755),
    .SCE(net772),
    .SET_B(net780),
    .Q(net595),
    .Q_N(net594));
 sky130_fd_sc_hd__a2111o_1 c733 (.A1(clknet_1_1__leaf_net556),
    .A2(clknet_1_1__leaf_net590),
    .B1(net549),
    .C1(net490),
    .D1(clknet_1_1__leaf_net755),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net578),
    .A1(net470),
    .A2(net565),
    .A3(net594),
    .S0(net947),
    .S1(clknet_1_0__leaf_net698),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net949),
    .A1(net575),
    .A2(clknet_1_1__leaf_net591),
    .A3(net470),
    .S0(net102),
    .S1(net947),
    .X(net598));
 sky130_fd_sc_hd__or4bb_1 c736 (.A(net934),
    .B(clknet_1_1__leaf_net556),
    .C_N(net594),
    .D_N(clknet_1_1__leaf_net699),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net817),
    .A1(clknet_1_1__leaf_net587),
    .A2(net339),
    .A3(net930),
    .S0(clknet_1_1__leaf_net755),
    .S1(net782),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net103),
    .A1(net339),
    .A2(net594),
    .A3(net780),
    .S0(net781),
    .S1(net783),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net473),
    .A1(net595),
    .A2(net549),
    .A3(net470),
    .S0(net947),
    .S1(net780),
    .X(net602));
 sky130_fd_sc_hd__a2111o_1 c74 (.A1(net5),
    .A2(net809),
    .B1(net7),
    .C1(net4),
    .D1(net951),
    .X(net11));
 sky130_fd_sc_hd__sdfbbp_1 c740 (.CLK(clknet_4_15_0_clk),
    .D(net941),
    .RESET_B(net565),
    .SCD(net470),
    .SCE(net595),
    .SET_B(net781),
    .Q(net603));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net533),
    .A1(net603),
    .A2(net472),
    .A3(net551),
    .S0(net781),
    .S1(net783),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_0__leaf_net590),
    .A1(net596),
    .A2(net533),
    .A3(net929),
    .S0(net779),
    .S1(net781),
    .X(net605));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(clknet_1_1__leaf_net591),
    .A2(net599),
    .B1(net70),
    .C1(net522),
    .D1(net783),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_0__leaf_net587),
    .A1(clknet_1_0__leaf_net591),
    .A2(net549),
    .A3(net938),
    .S0(net783),
    .S1(net785),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net938),
    .A1(net466),
    .A2(net490),
    .A3(net784),
    .S0(net785),
    .S1(net787),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net526),
    .A1(net601),
    .A2(clknet_1_0__leaf_net587),
    .A3(clknet_1_0__leaf_net591),
    .S0(net581),
    .S1(net786),
    .X(net609));
 sky130_fd_sc_hd__a2111o_1 c747 (.A1(net608),
    .A2(net595),
    .B1(clknet_1_1__leaf_net698),
    .C1(net779),
    .D1(net783),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net595),
    .A1(net947),
    .A2(net522),
    .A3(net574),
    .S0(clknet_1_1__leaf_net755),
    .S1(net766),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net522),
    .A1(net575),
    .A2(net930),
    .A3(net595),
    .S0(clknet_1_1__leaf_net517),
    .S1(net947),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c75 (.A0(net4),
    .A1(net880),
    .A2(net10),
    .A3(net7),
    .S0(net950),
    .S1(net16),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net611),
    .A1(net610),
    .A2(net929),
    .A3(net869),
    .S0(net595),
    .S1(net759),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net365),
    .A1(net490),
    .A2(net546),
    .A3(net869),
    .S0(net594),
    .S1(net766),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net614),
    .A1(net490),
    .A2(net365),
    .A3(net835),
    .S0(net574),
    .S1(net930),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net933),
    .A1(net489),
    .A2(net365),
    .A3(net818),
    .S0(net929),
    .S1(net766),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net604),
    .A1(net546),
    .A2(net930),
    .A3(net525),
    .S0(net594),
    .S1(net760),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net525),
    .A1(net612),
    .A2(net947),
    .A3(net930),
    .S0(net490),
    .S1(clknet_1_1__leaf_net755),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net930),
    .A1(net522),
    .A2(net546),
    .A3(net614),
    .S0(net759),
    .S1(net788),
    .X(net619));
 sky130_fd_sc_hd__a2111o_1 c757 (.A1(net619),
    .A2(net546),
    .B1(clknet_1_0__leaf_net517),
    .C1(net930),
    .D1(clknet_1_1__leaf_net756),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net411),
    .A1(net835),
    .A2(net522),
    .A3(clknet_1_0__leaf_net517),
    .S0(net760),
    .S1(net766),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net615),
    .A1(clknet_1_1__leaf_net621),
    .A2(net931),
    .A3(net594),
    .S0(net711),
    .S1(net766),
    .X(net622));
 sky130_fd_sc_hd__a2111o_1 c76 (.A1(net10),
    .A2(net23),
    .B1(net854),
    .C1(net6),
    .D1(net16),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(clknet_1_1__leaf_net517),
    .A1(net575),
    .A2(clknet_1_1__leaf_net621),
    .A3(net490),
    .S0(net696),
    .S1(net705),
    .X(net623));
 sky130_fd_sc_hd__a2111o_1 c761 (.A1(clknet_1_0__leaf_net621),
    .A2(net617),
    .B1(net623),
    .C1(net575),
    .D1(net930),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net606),
    .A1(net575),
    .A2(clknet_1_0__leaf_net621),
    .A3(net365),
    .S0(net704),
    .S1(net789),
    .X(net625));
 sky130_fd_sc_hd__and2_4 c77 (.A(net862),
    .B(net847),
    .X(net14));
 sky130_fd_sc_hd__and2_4 c78 (.A(net809),
    .B(net821),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c79 (.A(net839),
    .B(net15),
    .X(net16));
 sky130_fd_sc_hd__and2_4 c80 (.A(net809),
    .B(net854),
    .X(net17));
 sky130_fd_sc_hd__and2_2 c81 (.A(net835),
    .B(net855),
    .X(net918));
 sky130_fd_sc_hd__and2_2 c82 (.A(net857),
    .B(net850),
    .X(net18));
 sky130_fd_sc_hd__or4bb_4 c83 (.A(net15),
    .B(net951),
    .C_N(net819),
    .D_N(net950),
    .X(net19));
 sky130_fd_sc_hd__and3_4 c84 (.A(net19),
    .B(net950),
    .C(net823),
    .X(net20));
 sky130_fd_sc_hd__and2_0 c85 (.A(net818),
    .B(net20),
    .X(net21));
 sky130_fd_sc_hd__or4bb_2 c86 (.A(net853),
    .B(net20),
    .C_N(net15),
    .D_N(net844),
    .X(net22));
 sky130_fd_sc_hd__and2_1 c87 (.A(net835),
    .B(net851),
    .X(net23));
 sky130_fd_sc_hd__and3_1 c88 (.A(net9),
    .B(net3),
    .C(net862),
    .X(net24));
 sky130_fd_sc_hd__and2_4 c89 (.A(net24),
    .B(net8),
    .X(net25));
 sky130_fd_sc_hd__and2_1 c90 (.A(net812),
    .B(net958),
    .X(net26));
 sky130_fd_sc_hd__and2_2 c91 (.A(net844),
    .B(net836),
    .X(net27));
 sky130_fd_sc_hd__and2_1 c92 (.A(net3),
    .B(net27),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c93 (.A(net28),
    .B(net27),
    .X(net29));
 sky130_fd_sc_hd__and2_0 c94 (.A(net849),
    .B(net9),
    .X(net30));
 sky130_fd_sc_hd__and2_1 c95 (.A(net27),
    .B(net29),
    .X(net31));
 sky130_fd_sc_hd__and2_0 c96 (.A(net11),
    .B(net27),
    .X(net32));
 sky130_fd_sc_hd__and2_1 c97 (.A(net30),
    .B(net11),
    .X(net33));
 sky130_fd_sc_hd__and2_4 c98 (.A(net21),
    .B(net31),
    .X(net875));
 sky130_fd_sc_hd__and2_1 c99 (.A(net855),
    .B(net831),
    .X(net34));
 sky130_fd_sc_hd__or4bb_1 merge763 (.A(net315),
    .B(net198),
    .C_N(net952),
    .D_N(net703),
    .X(net626));
 sky130_fd_sc_hd__sdfbbn_1 merge764 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net870),
    .RESET_B(net189),
    .SCE(net243),
    .SET_B(net674),
    .Q(net340),
    .Q_N(net627));
 sky130_fd_sc_hd__clkbuf_1 merge765 (.A(net795),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 merge766 (.A0(net364),
    .A1(net367),
    .A2(net365),
    .A3(net927),
    .S0(net679),
    .S1(net722),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net445),
    .A1(net872),
    .A2(net437),
    .A3(net425),
    .S0(net453),
    .S1(net728),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 merge768 (.A0(net334),
    .A1(net929),
    .A2(net944),
    .A3(net310),
    .S0(net416),
    .S1(net433),
    .X(net632));
 sky130_fd_sc_hd__or4bb_1 merge769 (.A(net423),
    .B(net519),
    .C_N(net406),
    .D_N(net746),
    .X(net633));
 sky130_fd_sc_hd__a2111o_1 merge770 (.A1(net296),
    .A2(net198),
    .B1(clknet_1_1__leaf_net302),
    .C1(net203),
    .D1(net952),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 merge771 (.A0(net79),
    .A1(net205),
    .A2(net225),
    .A3(net221),
    .S0(net224),
    .S1(net67),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 merge772 (.A0(net105),
    .A1(net111),
    .A2(net850),
    .A3(net135),
    .S0(net131),
    .S1(net843),
    .X(net636));
 sky130_fd_sc_hd__sedfxbp_1 merge773 (.CLK(clknet_4_4_0_clk),
    .D(net127),
    .DE(net239),
    .SCD(net18),
    .SCE(clknet_1_1__leaf_net246),
    .Q(net638),
    .Q_N(net637));
 sky130_fd_sc_hd__or4bb_1 merge774 (.A(net860),
    .B(net203),
    .C_N(net406),
    .D_N(net66),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net26),
    .A1(net239),
    .A2(net821),
    .A3(clknet_1_0__leaf_net274),
    .S0(net3),
    .S1(net908),
    .X(net640));
 sky130_fd_sc_hd__a2111o_1 merge776 (.A1(net151),
    .A2(net156),
    .B1(net999),
    .C1(net957),
    .D1(net141),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net98),
    .A1(net104),
    .A2(net105),
    .A3(net67),
    .S0(net837),
    .S1(net118),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net426),
    .A1(net938),
    .A2(net933),
    .A3(net422),
    .S0(net332),
    .S1(net534),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 merge779 (.A0(net364),
    .A1(net327),
    .A2(net948),
    .A3(net453),
    .S0(net449),
    .S1(net355),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net348),
    .A1(net929),
    .A2(net943),
    .A3(net330),
    .S0(clknet_1_1__leaf_net316),
    .S1(net326),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net22),
    .A1(net907),
    .A2(net932),
    .A3(net908),
    .S0(net228),
    .S1(net683),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(clknet_1_1__leaf_net541),
    .A1(net546),
    .A2(net403),
    .A3(net534),
    .S0(net538),
    .S1(net531),
    .X(net647));
 sky130_fd_sc_hd__a2111o_1 merge783 (.A1(net234),
    .A2(net205),
    .B1(net235),
    .C1(net76),
    .D1(net201),
    .X(net648));
 sky130_fd_sc_hd__or4bb_1 merge784 (.A(net407),
    .B(net306),
    .C_N(net423),
    .D_N(net746),
    .X(net649));
 sky130_fd_sc_hd__sdfbbn_1 merge785 (.CLK_N(clknet_4_10_0_clk),
    .D(net528),
    .RESET_B(net520),
    .SCD(net403),
    .SCE(net407),
    .SET_B(clknet_1_0__leaf_net870),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__sdfbbp_1 merge786 (.CLK(clknet_4_8_0_clk),
    .D(net203),
    .RESET_B(net406),
    .SCD(net405),
    .SCE(net410),
    .SET_B(net75),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net251),
    .A1(net882),
    .A2(net928),
    .A3(net275),
    .S0(net280),
    .S1(net681),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net198),
    .A1(net101),
    .A2(net319),
    .A3(clknet_1_0__leaf_net322),
    .S0(net324),
    .S1(clknet_1_0__leaf_net887),
    .X(net655));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net243),
    .A1(net960),
    .A2(net128),
    .A3(net252),
    .S0(clknet_1_1__leaf_net246),
    .S1(net729),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net272),
    .A1(net26),
    .A2(net276),
    .A3(net275),
    .S0(clknet_1_0__leaf_net274),
    .S1(net716),
    .X(net657));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net260),
    .A1(net843),
    .A2(net102),
    .A3(net254),
    .S0(net232),
    .S1(net928),
    .X(net658));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(clknet_1_0__leaf_net316),
    .A1(net330),
    .A2(clknet_1_0__leaf_net246),
    .A3(net18),
    .S0(net857),
    .S1(net703),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(clknet_1_1__leaf_net312),
    .A1(clknet_1_1__leaf_net322),
    .A2(clknet_1_0__leaf_net887),
    .A3(net211),
    .S0(net426),
    .S1(net548),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(clknet_1_1__leaf_net309),
    .A1(clknet_1_1__leaf_net305),
    .A2(net297),
    .A3(net542),
    .S0(clknet_1_0__leaf_net541),
    .S1(net429),
    .X(net661));
 sky130_fd_sc_hd__and2_0 merge795 (.A(net387),
    .B(net390),
    .X(net662));
 sky130_fd_sc_hd__and2_0 merge796 (.A(net170),
    .B(net175),
    .X(net663));
 sky130_fd_sc_hd__dfrbp_1 merge797 (.CLK(clknet_4_2_0_clk),
    .D(net626),
    .RESET_B(net655),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_6_0_clk),
    .D(net359),
    .RESET_B(net361),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__dfrtn_1 merge799 (.CLK_N(clknet_4_9_0_clk),
    .D(net440),
    .RESET_B(net439),
    .Q(net668));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net588),
    .B(net592),
    .X(net669));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_5_0_clk),
    .D(net58),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_2 merge802 (.CLK(clknet_4_2_0_clk),
    .D(net295),
    .RESET_B(net314),
    .Q(net670));
 sky130_fd_sc_hd__dfrtp_1 merge803 (.CLK(clknet_4_5_0_clk),
    .RESET_B(net159),
    .Q(net163));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net146),
    .B(net132),
    .X(net672));
 sky130_fd_sc_hd__dfsbp_1 merge805 (.CLK(clknet_4_3_0_clk),
    .D(net337),
    .Q(net342),
    .Q_N(net673));
 sky130_fd_sc_hd__dfsbp_1 merge806 (.CLK(clknet_4_6_0_clk),
    .D(net474),
    .SET_B(net478),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_4_13_0_clk),
    .D(net496),
    .SET_B(net497),
    .Q(net677));
 sky130_fd_sc_hd__dfstp_1 merge808 (.CLK(clknet_4_11_0_clk),
    .D(net569),
    .SET_B(net571),
    .Q(net678));
 sky130_fd_sc_hd__dfstp_1 merge809 (.CLK(clknet_4_1_0_clk),
    .D(net258),
    .SET_B(net264),
    .Q(net679));
 sky130_fd_sc_hd__and2_0 merge810 (.A(net227),
    .B(net635),
    .X(net680));
 sky130_fd_sc_hd__dlrbn_1 merge811 (.D(net268),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net283),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlrbn_1 merge812 (.D(net642),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net122),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__dlrbp_1 merge813 (.D(net523),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net633),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dlrbp_1 merge814 (.D(net639),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net649),
    .Q(net688),
    .Q_N(net687));
 sky130_fd_sc_hd__dlrtn_1 merge815 (.D(net290),
    .GATE_N(clknet_4_7_0_clk),
    .RESET_B(net291),
    .Q(net881));
 sky130_fd_sc_hd__and2_0 merge816 (.A(net625),
    .B(net613),
    .X(net689));
 sky130_fd_sc_hd__dlrtn_1 merge817 (.D(net452),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net459),
    .Q(net690));
 sky130_fd_sc_hd__dlrtn_1 merge818 (.D(net554),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net555),
    .Q(net691));
 sky130_fd_sc_hd__dlrtp_1 merge819 (.D(net233),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net237),
    .Q(net692));
 sky130_fd_sc_hd__dlrtp_1 merge820 (.D(net441),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net631),
    .Q(net693));
 sky130_fd_sc_hd__dlrtp_1 merge821 (.D(net636),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net641),
    .Q(net694));
 sky130_fd_sc_hd__edfxbp_1 merge822 (.CLK(clknet_4_12_0_clk),
    .D(net689),
    .DE(net498),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__and2_0 merge823 (.A(net176),
    .B(net182),
    .X(net697));
 sky130_fd_sc_hd__edfxtp_1 merge824 (.CLK(clknet_4_7_0_clk),
    .D(net185),
    .DE(net662),
    .Q(net903));
 sky130_fd_sc_hd__sdlclkp_1 merge825 (.CLK(clknet_4_14_0_clk),
    .GATE(net593),
    .SCE(net609),
    .GCLK(net698));
 sky130_fd_sc_hd__sdlclkp_2 merge826 (.CLK(clknet_4_14_0_clk),
    .GATE(net576),
    .SCE(net669),
    .GCLK(net699));
 sky130_fd_sc_hd__sdlclkp_4 merge827 (.CLK(clknet_4_1_0_clk),
    .GATE(net266),
    .SCE(net648),
    .GCLK(net909));
 sky130_fd_sc_hd__dfrbp_1 merge828 (.CLK(clknet_4_13_0_clk),
    .D(net398),
    .RESET_B(net396),
    .Q(net883),
    .Q_N(net700));
 sky130_fd_sc_hd__dfrbp_1 merge829 (.CLK(clknet_4_2_0_clk),
    .D(net632),
    .RESET_B(net634),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__dfrtn_1 merge830 (.CLK_N(clknet_4_0_0_clk),
    .D(net202),
    .RESET_B(net680),
    .Q(net703));
 sky130_fd_sc_hd__dfrtp_1 merge831 (.CLK(clknet_4_15_0_clk),
    .D(net493),
    .RESET_B(net624),
    .Q(net704));
 sky130_fd_sc_hd__dfrtp_1 merge832 (.CLK(clknet_4_15_0_clk),
    .D(net509),
    .RESET_B(net622),
    .Q(net705));
 sky130_fd_sc_hd__dfrtp_1 merge833 (.CLK(clknet_4_0_0_clk),
    .RESET_B(net114),
    .Q(net120));
 sky130_fd_sc_hd__dfsbp_1 merge834 (.CLK(clknet_4_13_0_clk),
    .D(net501),
    .SET_B(net502),
    .Q(net708),
    .Q_N(net707));
 sky130_fd_sc_hd__dfsbp_2 merge835 (.CLK(clknet_4_1_0_clk),
    .D(net124),
    .SET_B(net672),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dfstp_1 merge836 (.CLK(clknet_4_13_0_clk),
    .D(net511),
    .SET_B(net620),
    .Q(net711));
 sky130_fd_sc_hd__dfstp_1 merge837 (.CLK(clknet_4_5_0_clk),
    .D(net663),
    .SET_B(net697),
    .Q(net900));
 sky130_fd_sc_hd__dfstp_1 merge838 (.CLK(clknet_4_2_0_clk),
    .D(net661),
    .SET_B(net659),
    .Q(net712));
 sky130_fd_sc_hd__dfxbp_1 s839 (.CLK(clknet_4_4_0_clk),
    .D(net144),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfxbp_1 s840 (.CLK(clknet_4_7_0_clk),
    .D(net162),
    .Q(net895),
    .Q_N(net715));
 sky130_fd_sc_hd__dfxtp_2 s841 (.CLK(clknet_4_4_0_clk),
    .D(net164),
    .Q(net884));
 sky130_fd_sc_hd__dfxtp_1 s842 (.CLK(clknet_4_5_0_clk),
    .D(net166),
    .Q(net716));
 sky130_fd_sc_hd__dfxtp_1 s843 (.CLK(clknet_4_5_0_clk),
    .D(net184),
    .Q(net901));
 sky130_fd_sc_hd__dlclkp_1 s844 (.CLK(clknet_4_4_0_clk),
    .GATE(net242),
    .GCLK(net717));
 sky130_fd_sc_hd__dlclkp_2 s845 (.CLK(clknet_4_1_0_clk),
    .GATE(net244),
    .GCLK(net718));
 sky130_fd_sc_hd__dlclkp_4 s846 (.CLK(clknet_4_1_0_clk),
    .GATE(net247),
    .GCLK(net719));
 sky130_fd_sc_hd__dlxbn_1 s847 (.D(net248),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlxbn_1 s848 (.D(net267),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dlxbp_1 s849 (.D(net278),
    .GATE(clknet_4_5_0_clk),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dlxtn_1 s850 (.D(net288),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net896));
 sky130_fd_sc_hd__dlxtn_1 s851 (.D(net289),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dlxtn_1 s852 (.D(net344),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net726));
 sky130_fd_sc_hd__dlxtp_1 s853 (.D(net350),
    .GATE(clknet_4_2_0_clk),
    .Q(net727));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s854 (.D(net351),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net728));
 sky130_fd_sc_hd__dfxbp_1 s855 (.CLK(clknet_4_6_0_clk),
    .D(net354),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dfxbp_1 s856 (.CLK(clknet_4_3_0_clk),
    .D(net357),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__dfxtp_1 s857 (.CLK(clknet_4_6_0_clk),
    .D(net374),
    .Q(net733));
 sky130_fd_sc_hd__dfxtp_1 s858 (.CLK(clknet_4_6_0_clk),
    .D(net375),
    .Q(net734));
 sky130_fd_sc_hd__dfxtp_1 s859 (.CLK(clknet_4_7_0_clk),
    .D(net379),
    .Q(net735));
 sky130_fd_sc_hd__dlclkp_1 s860 (.CLK(clknet_4_6_0_clk),
    .GATE(net380),
    .GCLK(net736));
 sky130_fd_sc_hd__dlclkp_2 s861 (.CLK(clknet_4_7_0_clk),
    .GATE(net382),
    .GCLK(net897));
 sky130_fd_sc_hd__dlclkp_4 s862 (.CLK(clknet_4_7_0_clk),
    .GATE(net384),
    .GCLK(net737));
 sky130_fd_sc_hd__dlxbn_1 s863 (.D(net385),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net739),
    .Q_N(net738));
 sky130_fd_sc_hd__dlxbn_1 s864 (.D(net386),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__dlxbp_1 s865 (.D(net388),
    .GATE(clknet_4_7_0_clk),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__dlxtn_1 s866 (.D(net389),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net891));
 sky130_fd_sc_hd__dlxtn_2 s867 (.D(net391),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net744));
 sky130_fd_sc_hd__dlxtn_2 s868 (.D(net420),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net745));
 sky130_fd_sc_hd__dlxtp_1 s869 (.D(net421),
    .GATE(clknet_4_8_0_clk),
    .Q(net746));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s870 (.D(net436),
    .SLEEP_B(clknet_4_9_0_clk),
    .Q(net747));
 sky130_fd_sc_hd__dfxbp_1 s871 (.CLK(clknet_4_12_0_clk),
    .D(net469),
    .Q(net749),
    .Q_N(net748));
 sky130_fd_sc_hd__dfxbp_1 s872 (.CLK(clknet_4_14_0_clk),
    .D(net471),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__dfxtp_1 s873 (.CLK(clknet_4_12_0_clk),
    .D(net483),
    .Q(net752));
 sky130_fd_sc_hd__dfxtp_1 s874 (.CLK(clknet_4_12_0_clk),
    .D(net484),
    .Q(net753));
 sky130_fd_sc_hd__dfxtp_1 s875 (.CLK(clknet_4_12_0_clk),
    .D(net485),
    .Q(net754));
 sky130_fd_sc_hd__dlclkp_1 s876 (.CLK(clknet_4_15_0_clk),
    .GATE(net495),
    .GCLK(net755));
 sky130_fd_sc_hd__dlclkp_2 s877 (.CLK(clknet_4_13_0_clk),
    .GATE(net499),
    .GCLK(net756));
 sky130_fd_sc_hd__dlclkp_4 s878 (.CLK(clknet_4_13_0_clk),
    .GATE(net500),
    .GCLK(net757));
 sky130_fd_sc_hd__dlxbn_1 s879 (.D(net504),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net758));
 sky130_fd_sc_hd__dlxbn_1 s880 (.D(net505),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dlxbp_1 s881 (.D(net506),
    .GATE(clknet_4_13_0_clk),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__dlxtn_2 s882 (.D(net507),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net877));
 sky130_fd_sc_hd__dlxtn_1 s883 (.D(net508),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net763));
 sky130_fd_sc_hd__dlxtn_1 s884 (.D(net512),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net764));
 sky130_fd_sc_hd__dlxtp_1 s885 (.D(net514),
    .GATE(clknet_4_13_0_clk),
    .Q(net765));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s886 (.D(net515),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net766));
 sky130_fd_sc_hd__dfxbp_1 s887 (.CLK(clknet_4_13_0_clk),
    .D(net516),
    .Q(net767));
 sky130_fd_sc_hd__dfxbp_1 s888 (.CLK(clknet_4_10_0_clk),
    .D(net535),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__dfxtp_2 s889 (.CLK(clknet_4_11_0_clk),
    .D(net558),
    .Q(net770));
 sky130_fd_sc_hd__dfxtp_1 s890 (.CLK(clknet_4_11_0_clk),
    .D(net562),
    .Q(net771));
 sky130_fd_sc_hd__dfxtp_1 s891 (.CLK(clknet_4_14_0_clk),
    .D(net579),
    .Q(net772));
 sky130_fd_sc_hd__dlclkp_1 s892 (.CLK(clknet_4_11_0_clk),
    .GATE(net580),
    .GCLK(net773));
 sky130_fd_sc_hd__dlclkp_2 s893 (.CLK(clknet_4_11_0_clk),
    .GATE(net582),
    .GCLK(net774));
 sky130_fd_sc_hd__dlclkp_4 s894 (.CLK(clknet_4_11_0_clk),
    .GATE(net584),
    .GCLK(net775));
 sky130_fd_sc_hd__dlxbn_1 s895 (.D(net585),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net777),
    .Q_N(net776));
 sky130_fd_sc_hd__dlxbn_1 s896 (.D(net586),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net778));
 sky130_fd_sc_hd__dlxbp_1 s897 (.D(net589),
    .GATE(clknet_4_14_0_clk),
    .Q(net780),
    .Q_N(net779));
 sky130_fd_sc_hd__dlxtn_1 s898 (.D(net597),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net781));
 sky130_fd_sc_hd__dlxtn_1 s899 (.D(net598),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net782));
 sky130_fd_sc_hd__dlxtn_1 s900 (.D(net600),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net783));
 sky130_fd_sc_hd__dlxtp_1 s901 (.D(net602),
    .GATE(clknet_4_14_0_clk),
    .Q(net784));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s902 (.D(net605),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net785));
 sky130_fd_sc_hd__dfxbp_1 s903 (.CLK(clknet_4_14_0_clk),
    .D(net607),
    .Q(net787),
    .Q_N(net786));
 sky130_fd_sc_hd__dfxbp_1 s904 (.CLK(clknet_4_12_0_clk),
    .D(net616),
    .Q(net788));
 sky130_fd_sc_hd__dfxtp_1 s905 (.CLK(clknet_4_15_0_clk),
    .D(net618),
    .Q(net789));
 sky130_fd_sc_hd__dfxtp_1 s906 (.CLK(clknet_4_3_0_clk),
    .D(net630),
    .Q(net790));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_4_0_clk),
    .D(net640),
    .Q(net791));
 sky130_fd_sc_hd__dlclkp_1 s908 (.CLK(clknet_4_10_0_clk),
    .GATE(net643),
    .GCLK(net792));
 sky130_fd_sc_hd__dlclkp_2 s909 (.CLK(clknet_4_12_0_clk),
    .GATE(net644),
    .GCLK(net793));
 sky130_fd_sc_hd__dlclkp_4 s910 (.CLK(clknet_4_2_0_clk),
    .GATE(net645),
    .GCLK(net794));
 sky130_fd_sc_hd__dlxbn_1 s911 (.D(net646),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net796),
    .Q_N(net795));
 sky130_fd_sc_hd__dlxbn_1 s912 (.D(net647),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net798),
    .Q_N(net797));
 sky130_fd_sc_hd__dlxbp_1 s913 (.D(net654),
    .GATE(clknet_4_4_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxtn_1 s914 (.D(net656),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net801));
 sky130_fd_sc_hd__dlxtn_1 s915 (.D(net657),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net802));
 sky130_fd_sc_hd__dlxtn_1 s916 (.D(net658),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net803));
 sky130_fd_sc_hd__dlxtp_1 s917 (.D(net660),
    .GATE(clknet_4_10_0_clk),
    .Q(net804));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net628));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net805));
 sky130_fd_sc_hd__buf_2 input3 (.A(in10),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in11),
    .X(net807));
 sky130_fd_sc_hd__buf_4 input5 (.A(in12),
    .X(net808));
 sky130_fd_sc_hd__buf_12 input6 (.A(in13),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(in15),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in17),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net814));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net815));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net816));
 sky130_fd_sc_hd__buf_4 input14 (.A(in20),
    .X(net817));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net818));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net820));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net822));
 sky130_fd_sc_hd__buf_1 input20 (.A(in26),
    .X(net823));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(in27),
    .X(net824));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net826));
 sky130_fd_sc_hd__buf_1 input24 (.A(in3),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input27 (.A(in32),
    .X(net830));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(in34),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in35),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in38),
    .X(net836));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(in40),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(in42),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(in43),
    .X(net842));
 sky130_fd_sc_hd__buf_4 input40 (.A(in44),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(in45),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input46 (.A(in5),
    .X(net849));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(in50),
    .X(net850));
 sky130_fd_sc_hd__buf_2 input48 (.A(in51),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net854));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net855));
 sky130_fd_sc_hd__buf_2 input53 (.A(in56),
    .X(net856));
 sky130_fd_sc_hd__buf_2 input54 (.A(in57),
    .X(net857));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(in58),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in59),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(in6),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in60),
    .X(net861));
 sky130_fd_sc_hd__buf_6 input59 (.A(in61),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input60 (.A(in7),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input61 (.A(in8),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(in9),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net866),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net867),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net868),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output66 (.A(net869),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(clknet_1_0__leaf_net870),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net871),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net872),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output70 (.A(net873),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output71 (.A(net874),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net875),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net876),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output74 (.A(net877),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output75 (.A(net936),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net879),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net880),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net881),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net882),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net883),
    .X(out25));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net884),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net885),
    .X(out27));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net886),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(clknet_1_1__leaf_net887),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net955),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output86 (.A(net889),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net890),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net891),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net892),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net893),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net894),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net895),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net896),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(clknet_1_1__leaf_net897),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net898),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output96 (.A(net899),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net900),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net901),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net902),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net903),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net904),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net905),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net906),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net907),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output105 (.A(net908),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(clknet_1_0__leaf_net909),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output107 (.A(net910),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net911),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net912),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net913),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net914),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net915),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net916),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net917),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output115 (.A(net918),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output116 (.A(net919),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net920),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net921),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net922),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output120 (.A(net923),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output121 (.A(net924),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(clknet_1_1__leaf_net925),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output123 (.A(net926),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net879),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net253),
    .X(net928));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net899),
    .X(net929));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net931),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net458),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net261),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net199),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net339),
    .X(net934));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net878),
    .X(net937));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net869),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net195),
    .X(net939));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net113),
    .X(net940));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net551),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net926),
    .X(net942));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net434),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net946),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_2 fanout142 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(net411),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout144 (.A(net411),
    .X(net947));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net892),
    .X(net948));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net70),
    .X(net949));
 sky130_fd_sc_hd__buf_12 fanout147 (.A(net17),
    .X(net950));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net14),
    .X(net951));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net297),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net298),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net794 (.A(net794),
    .X(clknet_0_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net568 (.A(net568),
    .X(clknet_0_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_0__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net568 (.A(clknet_0_net568),
    .X(clknet_1_1__leaf_net568));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net774 (.A(net774),
    .X(clknet_0_net774));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net774 (.A(clknet_0_net774),
    .X(clknet_1_0__leaf_net774));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net774 (.A(clknet_0_net774),
    .X(clknet_1_1__leaf_net774));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net591 (.A(net591),
    .X(clknet_0_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_0__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_1__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net698 (.A(net698),
    .X(clknet_0_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_0__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net698 (.A(clknet_0_net698),
    .X(clknet_1_1__leaf_net698));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net590 (.A(net590),
    .X(clknet_0_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_0__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_1__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net775 (.A(net775),
    .X(clknet_0_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_0__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net775 (.A(clknet_0_net775),
    .X(clknet_1_1__leaf_net775));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net587 (.A(net587),
    .X(clknet_0_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_0__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_1__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net333 (.A(net333),
    .X(clknet_0_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_0__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net737 (.A(net737),
    .X(clknet_0_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_0__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_1__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net793 (.A(net793),
    .X(clknet_0_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_0__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_1__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net360 (.A(net360),
    .X(clknet_0_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_0__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net360 (.A(clknet_0_net360),
    .X(clknet_1_1__leaf_net360));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net792 (.A(net792),
    .X(clknet_0_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net792 (.A(clknet_0_net792),
    .X(clknet_1_0__leaf_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net792 (.A(clknet_0_net792),
    .X(clknet_1_1__leaf_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net773 (.A(net773),
    .X(clknet_0_net773));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net773 (.A(clknet_0_net773),
    .X(clknet_1_0__leaf_net773));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net773 (.A(clknet_0_net773),
    .X(clknet_1_1__leaf_net773));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net583 (.A(net583),
    .X(clknet_0_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_0__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_1__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net541 (.A(net541),
    .X(clknet_0_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_0__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net541 (.A(clknet_0_net541),
    .X(clknet_1_1__leaf_net541));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net757 (.A(net757),
    .X(clknet_0_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_0__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net757 (.A(clknet_0_net757),
    .X(clknet_1_1__leaf_net757));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net517 (.A(net517),
    .X(clknet_0_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_0__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net517 (.A(clknet_0_net517),
    .X(clknet_1_1__leaf_net517));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net621 (.A(net621),
    .X(clknet_0_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_0__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net621 (.A(clknet_0_net621),
    .X(clknet_1_1__leaf_net621));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net756 (.A(net756),
    .X(clknet_0_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_0__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net756 (.A(clknet_0_net756),
    .X(clknet_1_1__leaf_net756));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net755 (.A(net755),
    .X(clknet_0_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net755 (.A(clknet_0_net755),
    .X(clknet_1_0__leaf_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net755 (.A(clknet_0_net755),
    .X(clknet_1_1__leaf_net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net736 (.A(net736),
    .X(clknet_0_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_0__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_1__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net925 (.A(net925),
    .X(clknet_0_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_0__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net925 (.A(clknet_0_net925),
    .X(clknet_1_1__leaf_net925));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(net961),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net265 (.A(net265),
    .X(clknet_0_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_0__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net265 (.A(clknet_0_net265),
    .X(clknet_1_1__leaf_net265));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net909 (.A(net909),
    .X(clknet_0_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_0__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net909 (.A(clknet_0_net909),
    .X(clknet_1_1__leaf_net909));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net238 (.A(net238),
    .X(clknet_0_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_0__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net238 (.A(clknet_0_net238),
    .X(clknet_1_1__leaf_net238));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net246 (.A(net246),
    .X(clknet_0_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_0__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net246 (.A(clknet_0_net246),
    .X(clknet_1_1__leaf_net246));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net718 (.A(net718),
    .X(clknet_0_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net718 (.A(clknet_0_net718),
    .X(clknet_1_0__leaf_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net718 (.A(clknet_0_net718),
    .X(clknet_1_1__leaf_net718));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net206 (.A(net206),
    .X(clknet_0_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_0__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net206 (.A(clknet_0_net206),
    .X(clknet_1_1__leaf_net206));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net312 (.A(net312),
    .X(clknet_0_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_0__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_1__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net322 (.A(net322),
    .X(clknet_0_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net322 (.A(clknet_0_net322),
    .X(clknet_1_0__leaf_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net322 (.A(clknet_0_net322),
    .X(clknet_1_1__leaf_net322));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net870 (.A(net870),
    .X(clknet_0_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net870 (.A(clknet_0_net870),
    .X(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net870 (.A(clknet_0_net870),
    .X(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net309 (.A(net309),
    .X(clknet_0_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_0__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_1__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net305 (.A(net305),
    .X(clknet_0_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_0__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net305 (.A(clknet_0_net305),
    .X(clknet_1_1__leaf_net305));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net717 (.A(net717),
    .X(clknet_0_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_0__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net717 (.A(clknet_0_net717),
    .X(clknet_1_1__leaf_net717));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net274 (.A(net274),
    .X(clknet_0_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_0__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net274 (.A(clknet_0_net274),
    .X(clknet_1_1__leaf_net274));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net699 (.A(net699),
    .X(clknet_0_net699));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net699 (.A(clknet_0_net699),
    .X(clknet_1_0__leaf_net699));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net699 (.A(clknet_0_net699),
    .X(clknet_1_1__leaf_net699));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net888),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net954),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net955),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net9),
    .X(net957));
 sky130_fd_sc_hd__and3_1 clone5 (.A(net19),
    .B(net950),
    .C(net823),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net19),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_1 clone7 (.A(net17),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(clknet_0_net397),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net951),
    .X(net962));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer10 (.A(net962),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net963),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net963),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net965),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net747),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net734),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net714),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net750),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net735),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net713),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net435),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net404),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net340),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net682),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net890),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net480),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net728),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net690),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net726),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net465),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net179),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net373),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net754),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net764),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net733),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net790),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net548),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net882),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net675),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net430),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net281),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net444),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net743),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net694),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net884),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net548),
    .X(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SCE (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCD (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCD (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_SET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SET_B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_C_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_Q_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_SCD (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_Q (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_C_N (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SCD (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_C1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A3 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_C1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_C_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_C (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_Q (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_SCD (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SCE (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SET_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_Q_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_X (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_SCD (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_RESET_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_C_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_D_N (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_D_N (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_C_N (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCD (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCD (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_D_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_RESET_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_RESET_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_DE (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_D (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_C (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_RESET_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_SCE (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_SCE (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SET_B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Q_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_Q (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_C1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_D_N (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_DE (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net333_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SCE (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_Q (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_SCE (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_Q (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_RESET_B (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_X (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCD (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCE (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_B1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_Q (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_Q_N (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_Q (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_X (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C_N (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_C (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A1 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C_N (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_C (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SCD (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_D (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_SCD (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_D1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SET_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_C1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_RESET_B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_D1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_SCE (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_X (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_C (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold20_A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_C1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_SCE (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_Q (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_X (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SCD (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A3 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCD (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_Q_N (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_SCD (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_X (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_C1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_X (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_D1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_C_N (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_B1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_D_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_X (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_RESET_B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_X (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_X (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_RESET_B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_RESET_B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_RESET_B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_X (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_C1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_Q_N (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_C1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_D_N (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_D1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_Q (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_D1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_C (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_Q (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SET_B (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S0 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Q (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_D1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_Q (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_Q_N (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_Q (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_C (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_SET_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_C (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_S1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_Q (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_C_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_D1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_D1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_D_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_C1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_C_N (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_C_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_D_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SCD (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_RESET_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_C1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_D_N (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_SCE (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_C (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_D1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SCE (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_D_N (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_C1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCD (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_C1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_C (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_D1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCD (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCE (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_S0 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_Q (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_D_N (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_Q (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_S1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net887_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_Q (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_C (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A0 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_SCD (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_C_N (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_SET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_S1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_C (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_C (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_Q (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_C1 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_S0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_D_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_RESET_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_SCD (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_SCE (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_RESET_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_RESET_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_B1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D_N (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_SCD (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_C1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_D1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_D1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_D_N (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C1 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_C (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_SCE (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCE (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_SET_B (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S0 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_C (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_B1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SCD (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCE (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_D_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_C (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_C (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_D_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_C1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_D_N (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_D1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C_N (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C_N (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_C_N (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_D1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_D_N (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_C (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_C (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C_N (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_D (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_C1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SCE (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCD (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_SCD (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCE (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_D1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_SET_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_D_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C_N (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_C1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_D_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_D1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_C (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_D_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_C_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_D1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_D_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_D_N (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_C (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_C (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_C (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_SCE (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s855_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_SLEEP_B (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_RESET_B (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_SCD (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_RESET_B (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net333_X (.DIODE(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_RESET_B (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net887_X (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net870_A (.DIODE(clknet_0_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net870_A (.DIODE(clknet_0_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net870_X (.DIODE(clknet_0_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_SCE (.DIODE(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_SCE (.DIODE(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SET_B (.DIODE(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net870_X (.DIODE(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_SCE (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_D (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net870_X (.DIODE(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_C1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_X (.DIODE(net960));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net38),
    .X(net999));
 sky130_fd_sc_hd__and2_1 clone6 (.A(net39),
    .B(net37),
    .X(net1000));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
