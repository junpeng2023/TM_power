module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net624;
 wire net693;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net806;
 wire clknet_1_0__leaf_net806;
 wire clknet_1_1__leaf_net806;
 wire clknet_0_net622;
 wire clknet_1_0__leaf_net622;
 wire clknet_1_1__leaf_net622;
 wire clknet_0_net708;
 wire clknet_1_0__leaf_net708;
 wire clknet_1_1__leaf_net708;
 wire clknet_0_net892;
 wire clknet_1_0__leaf_net892;
 wire clknet_1_1__leaf_net892;
 wire clknet_0_net789;
 wire clknet_1_0__leaf_net789;
 wire clknet_1_1__leaf_net789;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net480;
 wire clknet_1_0__leaf_net480;
 wire clknet_1_1__leaf_net480;
 wire clknet_0_net482;
 wire clknet_1_0__leaf_net482;
 wire clknet_1_1__leaf_net482;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net477;
 wire clknet_1_0__leaf_net477;
 wire clknet_1_1__leaf_net477;
 wire clknet_0_net771;
 wire clknet_1_0__leaf_net771;
 wire clknet_1_1__leaf_net771;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net770;
 wire clknet_1_0__leaf_net770;
 wire clknet_1_1__leaf_net770;
 wire clknet_0_net507;
 wire clknet_1_0__leaf_net507;
 wire clknet_1_1__leaf_net507;
 wire clknet_0_net769;
 wire clknet_1_0__leaf_net769;
 wire clknet_1_1__leaf_net769;
 wire clknet_0_net754;
 wire clknet_1_0__leaf_net754;
 wire clknet_1_1__leaf_net754;
 wire clknet_0_net168;
 wire clknet_1_0__leaf_net168;
 wire clknet_1_1__leaf_net168;
 wire clknet_0_net753;
 wire clknet_1_0__leaf_net753;
 wire clknet_1_1__leaf_net753;
 wire clknet_0_net930;
 wire clknet_1_0__leaf_net930;
 wire clknet_1_1__leaf_net930;
 wire clknet_0_net154;
 wire clknet_1_0__leaf_net154;
 wire clknet_1_1__leaf_net154;
 wire clknet_0_net752;
 wire clknet_1_0__leaf_net752;
 wire clknet_1_1__leaf_net752;
 wire clknet_0_net887;
 wire clknet_1_0__leaf_net887;
 wire clknet_1_1__leaf_net887;
 wire clknet_0_net919;
 wire clknet_1_0__leaf_net919;
 wire clknet_1_1__leaf_net919;
 wire clknet_0_net889;
 wire clknet_1_0__leaf_net889;
 wire clknet_1_1__leaf_net889;
 wire clknet_0_net744;
 wire clknet_1_0__leaf_net744;
 wire clknet_1_1__leaf_net744;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net344;
 wire clknet_1_0__leaf_net344;
 wire clknet_1_1__leaf_net344;
 wire clknet_0_net359;
 wire clknet_1_0__leaf_net359;
 wire clknet_1_1__leaf_net359;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net373;
 wire clknet_1_0__leaf_net373;
 wire clknet_1_1__leaf_net373;
 wire clknet_0_net376;
 wire clknet_1_0__leaf_net376;
 wire clknet_1_1__leaf_net376;
 wire clknet_0_net710;
 wire clknet_1_0__leaf_net710;
 wire clknet_1_1__leaf_net710;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;

 sky130_fd_sc_hd__and3_4 c100 (.A(net876),
    .B(net14),
    .C(net32),
    .X(net37));
 sky130_fd_sc_hd__and3_1 c101 (.A(net25),
    .B(net959),
    .C(net37),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net34),
    .A1(net37),
    .A2(net918),
    .A3(net32),
    .S0(net28),
    .S1(net999),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net38),
    .A1(net32),
    .A2(net39),
    .A3(net28),
    .S0(net26),
    .S1(net33),
    .X(net40));
 sky130_fd_sc_hd__a2111o_4 c104 (.A1(net27),
    .A2(net983),
    .B1(net39),
    .C1(net959),
    .D1(net950),
    .X(net41));
 sky130_fd_sc_hd__or4bb_2 c105 (.A(net30),
    .B(net37),
    .C_N(net36),
    .D_N(net39),
    .X(net42));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net35),
    .A1(net34),
    .A2(net25),
    .A3(net38),
    .S0(net41),
    .S1(net39),
    .X(net43));
 sky130_fd_sc_hd__or4bb_1 c107 (.A(net33),
    .B(net42),
    .C_N(net37),
    .X(net44));
 sky130_fd_sc_hd__a2111o_2 c108 (.A1(net39),
    .A2(net38),
    .B1(net959),
    .C1(net22),
    .D1(net701),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net33),
    .A1(net42),
    .A2(net26),
    .A3(net832),
    .S0(net959),
    .S1(net701),
    .X(net46));
 sky130_fd_sc_hd__and3_4 c110 (.A(net879),
    .B(net918),
    .C(net22),
    .X(net47));
 sky130_fd_sc_hd__and2_1 c111 (.A(net854),
    .B(net47),
    .X(net48));
 sky130_fd_sc_hd__and2_0 c112 (.A(net22),
    .B(net26),
    .X(net49));
 sky130_fd_sc_hd__and3_1 c113 (.A(net49),
    .B(net976),
    .C(net48),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 c114 (.A0(net48),
    .A1(net41),
    .A2(net50),
    .A3(net47),
    .S0(net977),
    .S1(net1062),
    .X(net51));
 sky130_fd_sc_hd__and2_0 c115 (.A(net49),
    .B(net888),
    .X(net52));
 sky130_fd_sc_hd__and2_1 c116 (.A(net50),
    .B(net1066),
    .X(net921));
 sky130_fd_sc_hd__and3_1 c117 (.A(net950),
    .B(net876),
    .C(net52),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c118 (.A(net50),
    .B(net36),
    .X(net54));
 sky130_fd_sc_hd__sdfrbp_1 c119 (.CLK(clknet_4_10_0_clk),
    .D(net48),
    .RESET_B(net47),
    .SCD(net49),
    .SCE(net41),
    .Q(net56),
    .Q_N(net55));
 sky130_fd_sc_hd__mux4_1 c120 (.A0(net36),
    .A1(net54),
    .A2(net56),
    .A3(net47),
    .S0(net53),
    .S1(net879),
    .X(net57));
 sky130_fd_sc_hd__and2_1 c121 (.A(net861),
    .B(net748),
    .X(net928));
 sky130_fd_sc_hd__and3_1 c122 (.A(net56),
    .B(net928),
    .C(net37),
    .X(net58));
 sky130_fd_sc_hd__buf_1 c123 (.A(net727),
    .X(net933));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net53),
    .A1(net48),
    .A2(net58),
    .A3(net37),
    .S0(net47),
    .S1(net1064),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 c125 (.A(net822),
    .X(net60));
 sky130_fd_sc_hd__and3_1 c126 (.A(net26),
    .B(net48),
    .C(net1067),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 c127 (.A(net727),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net56),
    .A1(net61),
    .A2(net48),
    .A3(net47),
    .S0(net50),
    .S1(net746),
    .X(net923));
 sky130_fd_sc_hd__or4bb_1 c129 (.A(net52),
    .B(net47),
    .C_N(net933),
    .D_N(net1029),
    .X(net936));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net876),
    .A1(net61),
    .A2(net936),
    .A3(net1038),
    .S0(net921),
    .S1(net1029),
    .X(net63));
 sky130_fd_sc_hd__mux4_2 c131 (.A0(net47),
    .A1(net936),
    .A2(net928),
    .A3(net847),
    .S0(net888),
    .S1(net749),
    .X(net64));
 sky130_fd_sc_hd__and3_4 c132 (.A(net882),
    .B(net828),
    .C(net835),
    .X(net65));
 sky130_fd_sc_hd__and3_4 c133 (.A(net835),
    .B(net832),
    .C(net878),
    .X(net66));
 sky130_fd_sc_hd__and3_4 c134 (.A(net66),
    .B(net65),
    .C(net826),
    .X(net67));
 sky130_fd_sc_hd__and3_2 c135 (.A(net693),
    .B(net65),
    .C(net827),
    .X(net68));
 sky130_fd_sc_hd__and3_4 c136 (.A(net67),
    .B(net881),
    .C(net832),
    .X(net69));
 sky130_fd_sc_hd__and3_2 c137 (.A(net65),
    .B(net826),
    .C(net833),
    .X(net70));
 sky130_fd_sc_hd__and3_4 c138 (.A(net69),
    .B(net66),
    .C(net70),
    .X(net894));
 sky130_fd_sc_hd__and3_1 c139 (.A(net70),
    .B(net833),
    .C(net882),
    .X(net71));
 sky130_fd_sc_hd__a2111o_2 c140 (.A1(net70),
    .A2(net71),
    .B1(net66),
    .C1(net69),
    .D1(net67),
    .X(net72));
 sky130_fd_sc_hd__and3_2 c141 (.A(net964),
    .B(net69),
    .C(net71),
    .X(net73));
 sky130_fd_sc_hd__and3_1 c142 (.A(net881),
    .B(net73),
    .C(net878),
    .X(net74));
 sky130_fd_sc_hd__mux4_2 c143 (.A0(net824),
    .A1(net826),
    .A2(net70),
    .A3(net68),
    .S0(net964),
    .S1(net624),
    .X(net75));
 sky130_fd_sc_hd__and3_2 c144 (.A(net73),
    .B(net974),
    .C(net72),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net65),
    .A1(net72),
    .A2(net74),
    .A3(net70),
    .S0(net836),
    .S1(net75),
    .X(net77));
 sky130_fd_sc_hd__and3_2 c146 (.A(net831),
    .B(net74),
    .C(net69),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c147 (.A(net827),
    .B(net74),
    .C(net824),
    .X(net79));
 sky130_fd_sc_hd__and3_1 c148 (.A(net66),
    .B(net73),
    .C(net881),
    .X(net80));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net833),
    .A1(net80),
    .A2(net79),
    .A3(net75),
    .S0(net832),
    .S1(net828),
    .X(net81));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net78),
    .A1(net81),
    .A2(net824),
    .A3(net77),
    .S0(net70),
    .S1(net867),
    .X(net82));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net74),
    .A1(net829),
    .A2(net82),
    .A3(net81),
    .S0(net964),
    .S1(net73),
    .X(net83));
 sky130_fd_sc_hd__and3_4 c152 (.A(net83),
    .B(net81),
    .C(net72),
    .X(net84));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net845),
    .A1(net83),
    .A2(net80),
    .A3(net84),
    .S0(net992),
    .S1(net82),
    .X(net85));
 sky130_fd_sc_hd__and2_2 c154 (.A(net843),
    .B(net883),
    .X(net86));
 sky130_fd_sc_hd__and2_4 c155 (.A(net75),
    .B(net853),
    .X(net885));
 sky130_fd_sc_hd__and3_1 c156 (.A(net846),
    .B(net76),
    .C(net84),
    .X(net87));
 sky130_fd_sc_hd__and3_1 c157 (.A(net86),
    .B(net962),
    .C(net846),
    .X(net88));
 sky130_fd_sc_hd__and2_4 c158 (.A(net838),
    .B(net87),
    .X(net89));
 sky130_fd_sc_hd__and2_0 c159 (.A(net857),
    .B(net84),
    .X(net90));
 sky130_fd_sc_hd__and2_1 c160 (.A(net853),
    .B(net962),
    .X(net91));
 sky130_fd_sc_hd__and2_4 c161 (.A(net855),
    .B(net838),
    .X(net92));
 sky130_fd_sc_hd__and2_2 c162 (.A(net88),
    .B(net91),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c163 (.A(net850),
    .B(net851),
    .X(net94));
 sky130_fd_sc_hd__a2111o_1 c164 (.A1(net860),
    .A2(net92),
    .B1(net91),
    .C1(net93),
    .D1(net84),
    .X(net95));
 sky130_fd_sc_hd__and2_2 c165 (.A(net93),
    .B(net95),
    .X(net96));
 sky130_fd_sc_hd__or4bb_4 c166 (.A(net91),
    .B(net90),
    .C_N(net852),
    .D_N(net859),
    .X(net97));
 sky130_fd_sc_hd__and2_2 c167 (.A(net844),
    .B(net95),
    .X(net98));
 sky130_fd_sc_hd__or4bb_1 c168 (.A(net856),
    .B(net87),
    .C_N(net93),
    .D_N(net987),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c169 (.A0(net99),
    .A1(net856),
    .A2(net93),
    .A3(net84),
    .S0(net89),
    .S1(net94),
    .X(net100));
 sky130_fd_sc_hd__and2_2 c170 (.A(net97),
    .B(net87),
    .X(net101));
 sky130_fd_sc_hd__and2_1 c171 (.A(net87),
    .B(net96),
    .X(net102));
 sky130_fd_sc_hd__and2_1 c172 (.A(net98),
    .B(net102),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net954),
    .A1(net843),
    .A2(net103),
    .A3(net97),
    .S0(net87),
    .S1(net98),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net99),
    .A1(net88),
    .A2(net89),
    .A3(net98),
    .S0(net954),
    .S1(net688),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net90),
    .A1(net837),
    .A2(net860),
    .A3(net842),
    .S0(net105),
    .X(net106));
 sky130_fd_sc_hd__and3_1 c176 (.A(net68),
    .B(net93),
    .C(net688),
    .X(net107));
 sky130_fd_sc_hd__and3_1 c177 (.A(net100),
    .B(net837),
    .C(net878),
    .X(net108));
 sky130_fd_sc_hd__buf_1 c178 (.A(net722),
    .X(net109));
 sky130_fd_sc_hd__and3_1 c179 (.A(net851),
    .B(net862),
    .C(net3),
    .X(net110));
 sky130_fd_sc_hd__and3_1 c180 (.A(net880),
    .B(net872),
    .C(net825),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c181 (.A(net111),
    .B(net837),
    .C(net863),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 c182 (.A(net722),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c183 (.A(net93),
    .B(net109),
    .C(net86),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 c184 (.A(net723),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c185 (.A(net3),
    .B(net113),
    .C(net873),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c186 (.A(net107),
    .B(net871),
    .C(net880),
    .X(net117));
 sky130_fd_sc_hd__a2111o_1 c187 (.A1(net115),
    .A2(net851),
    .B1(net966),
    .C1(net879),
    .D1(net109),
    .X(net118));
 sky130_fd_sc_hd__and3_1 c188 (.A(net117),
    .B(net965),
    .C(net109),
    .X(net119));
 sky130_fd_sc_hd__or4bb_4 c189 (.A(net875),
    .B(net873),
    .C_N(net119),
    .D_N(net965),
    .X(net120));
 sky130_fd_sc_hd__or4bb_1 c190 (.A(net119),
    .B(net120),
    .C_N(net109),
    .D_N(net965),
    .X(net121));
 sky130_fd_sc_hd__or4bb_1 c191 (.A(net109),
    .B(net100),
    .C_N(net111),
    .D_N(net965),
    .X(net122));
 sky130_fd_sc_hd__or4bb_4 c192 (.A(net121),
    .B(net76),
    .C_N(net965),
    .D_N(net873),
    .X(net123));
 sky130_fd_sc_hd__and3_1 c193 (.A(net117),
    .B(net965),
    .C(net953),
    .X(net124));
 sky130_fd_sc_hd__a2111o_4 c194 (.A1(net117),
    .A2(net110),
    .B1(net107),
    .C1(net93),
    .D1(net688),
    .X(net125));
 sky130_fd_sc_hd__a2111o_1 c195 (.A1(net112),
    .A2(net120),
    .B1(net965),
    .C1(net92),
    .D1(net688),
    .X(net126));
 sky130_fd_sc_hd__a2111o_1 c196 (.A1(net122),
    .A2(net125),
    .B1(net86),
    .C1(net112),
    .D1(net965),
    .X(net127));
 sky130_fd_sc_hd__sdfbbn_1 c197 (.CLK_N(clknet_4_2_0_clk),
    .D(net119),
    .RESET_B(net124),
    .SCD(net117),
    .SCE(net965),
    .SET_B(net723),
    .Q(net129),
    .Q_N(net128));
 sky130_fd_sc_hd__and3_1 c198 (.A(net842),
    .B(net125),
    .C(net69),
    .X(net130));
 sky130_fd_sc_hd__buf_1 c199 (.A(net737),
    .X(net131));
 sky130_fd_sc_hd__a2111o_1 c200 (.A1(net19),
    .A2(net998),
    .B1(net825),
    .C1(net17),
    .D1(net953),
    .X(net132));
 sky130_fd_sc_hd__sdfbbn_1 c201 (.CLK_N(clknet_4_2_0_clk),
    .D(net130),
    .RESET_B(net862),
    .SCD(net131),
    .SCE(net105),
    .SET_B(net965),
    .Q(net134),
    .Q_N(net133));
 sky130_fd_sc_hd__a2111o_4 c202 (.A1(net17),
    .A2(net113),
    .B1(net131),
    .C1(net125),
    .D1(net92),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 c203 (.A(net737),
    .X(net136));
 sky130_fd_sc_hd__and3_2 c204 (.A(net136),
    .B(net17),
    .C(net23),
    .X(net137));
 sky130_fd_sc_hd__and3_1 c205 (.A(net131),
    .B(net869),
    .C(net136),
    .X(net138));
 sky130_fd_sc_hd__a2111o_1 c206 (.A1(net132),
    .A2(net137),
    .B1(net832),
    .C1(net105),
    .D1(net134),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c207 (.A(net870),
    .B(net19),
    .C(net138),
    .X(net140));
 sky130_fd_sc_hd__a2111o_4 c208 (.A1(net137),
    .A2(net136),
    .B1(net128),
    .C1(net19),
    .D1(net135),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 c209 (.A(net730),
    .X(net142));
 sky130_fd_sc_hd__mux4_2 c210 (.A0(net142),
    .A1(net141),
    .A2(net134),
    .A3(net136),
    .S0(net138),
    .S1(net862),
    .X(net143));
 sky130_fd_sc_hd__a2111o_4 c211 (.A1(net143),
    .A2(net118),
    .B1(net130),
    .C1(net865),
    .D1(net128),
    .X(net920));
 sky130_fd_sc_hd__and3_4 c212 (.A(net140),
    .B(net143),
    .C(net141),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_4 c213 (.A(net737),
    .X(net144));
 sky130_fd_sc_hd__a2111o_1 c214 (.A1(net125),
    .A2(net143),
    .B1(net137),
    .C1(net23),
    .D1(net737),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(net138),
    .A1(net89),
    .A2(net979),
    .A3(net144),
    .S0(net145),
    .S1(net868),
    .X(net146));
 sky130_fd_sc_hd__a2111o_1 c216 (.A1(net852),
    .A2(net937),
    .B1(net847),
    .C1(net140),
    .D1(net138),
    .X(net147));
 sky130_fd_sc_hd__mux4_2 c217 (.A0(net138),
    .A1(net23),
    .A2(net141),
    .A3(net144),
    .S0(net136),
    .S1(net751),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net118),
    .A1(net143),
    .A2(net137),
    .A3(net148),
    .S0(net144),
    .S1(net751),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net149),
    .A1(net980),
    .A2(net96),
    .A3(net134),
    .S0(net737),
    .S1(net751),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 c220 (.A(net645),
    .X(net151));
 sky130_fd_sc_hd__and2_1 c221 (.A(net151),
    .B(net5),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c222 (.A0(net32),
    .A1(net148),
    .A2(net937),
    .A3(net33),
    .S0(net950),
    .S1(clknet_1_0__leaf_net752),
    .X(net153));
 sky130_fd_sc_hd__or4bb_1 c223 (.A(net869),
    .B(net5),
    .C_N(net967),
    .D_N(clknet_1_1__leaf_net752),
    .X(net887));
 sky130_fd_sc_hd__a2111o_1 c224 (.A1(net137),
    .A2(net1000),
    .B1(net25),
    .C1(net834),
    .D1(clknet_1_0__leaf_net753),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 c225 (.A(net645),
    .X(net155));
 sky130_fd_sc_hd__a2111o_1 c226 (.A1(net155),
    .A2(net874),
    .B1(net89),
    .C1(net37),
    .D1(clknet_1_0__leaf_net753),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net45),
    .A1(net36),
    .A2(net155),
    .A3(net69),
    .S0(net41),
    .S1(clknet_1_1__leaf_net753),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 c228 (.A(net823),
    .X(net158));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(net158),
    .A2(net148),
    .B1(net959),
    .C1(net41),
    .D1(clknet_1_1__leaf_net753),
    .X(net159));
 sky130_fd_sc_hd__or4bb_1 c230 (.A(net151),
    .B(net962),
    .C_N(clknet_1_0__leaf_net752),
    .D_N(clknet_1_0__leaf_net753),
    .X(net930));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net953),
    .A1(clknet_1_0__leaf_net930),
    .A2(net137),
    .A3(net155),
    .S0(net33),
    .S1(clknet_1_0__leaf_net752),
    .X(net160));
 sky130_fd_sc_hd__and2_1 c232 (.A(net152),
    .B(net743),
    .X(net161));
 sky130_fd_sc_hd__sdfbbp_1 c233 (.CLK(clknet_4_8_0_clk),
    .D(net1014),
    .RESET_B(net5),
    .SCD(clknet_1_0__leaf_net154),
    .SCE(net998),
    .SET_B(net41),
    .Q(net163),
    .Q_N(net162));
 sky130_fd_sc_hd__mux4_1 c234 (.A0(net42),
    .A1(net155),
    .A2(clknet_1_0__leaf_net154),
    .A3(clknet_1_1__leaf_net930),
    .S0(net979),
    .S1(net743),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 c235 (.A(net653),
    .X(net925));
 sky130_fd_sc_hd__and2_1 c236 (.A(net69),
    .B(net32),
    .X(net926));
 sky130_fd_sc_hd__buf_1 c237 (.A(net652),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net1001),
    .A1(net148),
    .A2(net162),
    .A3(net900),
    .S0(clknet_1_1__leaf_net753),
    .S1(clknet_1_1__leaf_net754),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net42),
    .A1(net925),
    .A2(net883),
    .A3(net155),
    .S0(net161),
    .S1(clknet_1_1__leaf_net754),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net163),
    .A1(net165),
    .A2(net925),
    .A3(net979),
    .S0(clknet_1_1__leaf_net753),
    .S1(clknet_1_0__leaf_net754),
    .X(net168));
 sky130_fd_sc_hd__buf_2 c241 (.A(net660),
    .X(net927));
 sky130_fd_sc_hd__and3_1 c242 (.A(net144),
    .B(net62),
    .C(net36),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_1 c243 (.A(net816),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_1 c244 (.A(net816),
    .X(net169));
 sky130_fd_sc_hd__and2_1 c245 (.A(net950),
    .B(net749),
    .X(net170));
 sky130_fd_sc_hd__buf_1 c246 (.A(net727),
    .X(net903));
 sky130_fd_sc_hd__and2_2 c247 (.A(net152),
    .B(net847),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 c248 (.A(net727),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net743),
    .X(net173));
 sky130_fd_sc_hd__and3_1 c250 (.A(net967),
    .B(net976),
    .C(net750),
    .X(net924));
 sky130_fd_sc_hd__and3_1 c251 (.A(net169),
    .B(net171),
    .C(net750),
    .X(net174));
 sky130_fd_sc_hd__and3_1 c252 (.A(net862),
    .B(net967),
    .C(net975),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net173),
    .A1(net41),
    .A2(net171),
    .A3(net967),
    .S0(net920),
    .S1(net749),
    .X(net176));
 sky130_fd_sc_hd__buf_1 c254 (.A(net743),
    .X(net177));
 sky130_fd_sc_hd__and3_4 c255 (.A(net64),
    .B(net37),
    .C(net757),
    .X(net911));
 sky130_fd_sc_hd__mux4_1 c256 (.A0(net165),
    .A1(net37),
    .A2(net911),
    .A3(net920),
    .S0(net171),
    .S1(net756),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 c257 (.A(net823),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_1 c258 (.A(net822),
    .X(net179));
 sky130_fd_sc_hd__a2111o_1 c259 (.A1(net174),
    .A2(net911),
    .B1(net152),
    .C1(clknet_1_1__leaf_net887),
    .D1(net757),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 c260 (.A(net659),
    .X(net902));
 sky130_fd_sc_hd__a2111o_1 c261 (.A1(net175),
    .A2(net170),
    .B1(net171),
    .C1(net911),
    .D1(net177),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net156),
    .A1(net171),
    .A2(net78),
    .A3(net726),
    .S0(net750),
    .S1(net755),
    .X(net910));
 sky130_fd_sc_hd__a2111o_1 c263 (.A1(net62),
    .A2(net165),
    .B1(net902),
    .C1(net883),
    .D1(net967),
    .X(net934));
 sky130_fd_sc_hd__and3_1 c264 (.A(net856),
    .B(net882),
    .C(net828),
    .X(net182));
 sky130_fd_sc_hd__and2_1 c265 (.A(net878),
    .B(net80),
    .X(net183));
 sky130_fd_sc_hd__and2_0 c266 (.A(net825),
    .B(net974),
    .X(net184));
 sky130_fd_sc_hd__and2_4 c267 (.A(net82),
    .B(net77),
    .X(net185));
 sky130_fd_sc_hd__and2_0 c268 (.A(net624),
    .B(net82),
    .X(net186));
 sky130_fd_sc_hd__and2_1 c269 (.A(net883),
    .B(net845),
    .X(net187));
 sky130_fd_sc_hd__and2_0 c270 (.A(net79),
    .B(net972),
    .X(net188));
 sky130_fd_sc_hd__and3_1 c271 (.A(net186),
    .B(net185),
    .C(net972),
    .X(net189));
 sky130_fd_sc_hd__and3_1 c272 (.A(net182),
    .B(net183),
    .C(net972),
    .X(net190));
 sky130_fd_sc_hd__and2_1 c273 (.A(net185),
    .B(net82),
    .X(net191));
 sky130_fd_sc_hd__and2_0 c274 (.A(net189),
    .B(net883),
    .X(net192));
 sky130_fd_sc_hd__and3_1 c275 (.A(net972),
    .B(net189),
    .C(net1011),
    .X(net193));
 sky130_fd_sc_hd__and2_0 c276 (.A(net193),
    .B(net76),
    .X(net194));
 sky130_fd_sc_hd__and2_2 c277 (.A(net80),
    .B(net67),
    .X(net195));
 sky130_fd_sc_hd__and3_1 c278 (.A(net189),
    .B(net835),
    .C(net972),
    .X(net196));
 sky130_fd_sc_hd__and2_1 c279 (.A(net182),
    .B(net972),
    .X(net197));
 sky130_fd_sc_hd__and3_2 c280 (.A(net194),
    .B(net79),
    .C(net972),
    .X(net938));
 sky130_fd_sc_hd__or4bb_4 c281 (.A(net196),
    .B(net952),
    .C_N(net867),
    .D_N(net972),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 c282 (.A(net729),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net192),
    .A1(net198),
    .A2(net199),
    .A3(net184),
    .S0(net829),
    .S1(net194),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net199),
    .A1(net198),
    .A2(net186),
    .A3(net952),
    .S0(net84),
    .S1(net829),
    .X(net201));
 sky130_fd_sc_hd__a2111o_4 c285 (.A1(net952),
    .A2(net882),
    .B1(net998),
    .C1(net972),
    .D1(net729),
    .X(net202));
 sky130_fd_sc_hd__and3_1 c286 (.A(net98),
    .B(net839),
    .C(net195),
    .X(net203));
 sky130_fd_sc_hd__and2_1 c287 (.A(net188),
    .B(net75),
    .X(net204));
 sky130_fd_sc_hd__and2_4 c288 (.A(net204),
    .B(net688),
    .X(net205));
 sky130_fd_sc_hd__and3_1 c289 (.A(net839),
    .B(net859),
    .C(net193),
    .X(net206));
 sky130_fd_sc_hd__and2_0 c290 (.A(net882),
    .B(net188),
    .X(net207));
 sky130_fd_sc_hd__and2_2 c291 (.A(net192),
    .B(net204),
    .X(net208));
 sky130_fd_sc_hd__buf_1 c292 (.A(net730),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c293 (.A(net207),
    .B(net183),
    .C(net190),
    .X(net210));
 sky130_fd_sc_hd__and3_1 c294 (.A(net203),
    .B(net206),
    .C(net210),
    .X(net211));
 sky130_fd_sc_hd__and2_1 c295 (.A(net102),
    .B(net205),
    .X(net212));
 sky130_fd_sc_hd__or4bb_1 c296 (.A(net188),
    .B(net212),
    .C_N(net103),
    .D_N(net954),
    .X(net213));
 sky130_fd_sc_hd__and3_1 c297 (.A(net210),
    .B(net193),
    .C(net688),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 c298 (.A(net728),
    .X(net215));
 sky130_fd_sc_hd__and2_0 c299 (.A(net849),
    .B(net207),
    .X(net216));
 sky130_fd_sc_hd__buf_1 c300 (.A(net728),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 c301 (.A(net729),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c302 (.A(net94),
    .B(net215),
    .C(net218),
    .X(net219));
 sky130_fd_sc_hd__and2_1 c303 (.A(net215),
    .B(net209),
    .X(net220));
 sky130_fd_sc_hd__and2_2 c304 (.A(net206),
    .B(net204),
    .X(net221));
 sky130_fd_sc_hd__or4bb_2 c305 (.A(net216),
    .B(net79),
    .C_N(net220),
    .D_N(net219),
    .X(net222));
 sky130_fd_sc_hd__and3_4 c306 (.A(net204),
    .B(net97),
    .C(net222),
    .X(net899));
 sky130_fd_sc_hd__mux4_2 c307 (.A0(net217),
    .A1(net215),
    .A2(net221),
    .A3(net839),
    .S0(net102),
    .S1(net195),
    .X(net223));
 sky130_fd_sc_hd__and2_0 c308 (.A(net95),
    .B(net197),
    .X(net224));
 sky130_fd_sc_hd__and3_2 c309 (.A(net837),
    .B(net962),
    .C(net95),
    .X(net225));
 sky130_fd_sc_hd__buf_1 c310 (.A(net686),
    .X(net226));
 sky130_fd_sc_hd__and3_2 c311 (.A(net865),
    .B(net113),
    .C(net688),
    .X(net227));
 sky130_fd_sc_hd__mux4_2 c312 (.A0(net879),
    .A1(net837),
    .A2(net113),
    .A3(net224),
    .S0(net958),
    .S1(net835),
    .X(net228));
 sky130_fd_sc_hd__and3_2 c313 (.A(net214),
    .B(net76),
    .C(net968),
    .X(net229));
 sky130_fd_sc_hd__buf_1 c314 (.A(net686),
    .X(net230));
 sky130_fd_sc_hd__and2_0 c315 (.A(net76),
    .B(net958),
    .X(net231));
 sky130_fd_sc_hd__and3_1 c316 (.A(net873),
    .B(net968),
    .C(net688),
    .X(net232));
 sky130_fd_sc_hd__and3_2 c317 (.A(net219),
    .B(net230),
    .C(net966),
    .X(net233));
 sky130_fd_sc_hd__and3_2 c318 (.A(net195),
    .B(net873),
    .C(net729),
    .X(net234));
 sky130_fd_sc_hd__and3_1 c319 (.A(net231),
    .B(net208),
    .C(net234),
    .X(net235));
 sky130_fd_sc_hd__and3_2 c320 (.A(net193),
    .B(net214),
    .C(net963),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 c321 (.A(net723),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 c322 (.A(net686),
    .X(net238));
 sky130_fd_sc_hd__mux4_2 c323 (.A0(net197),
    .A1(net226),
    .A2(net237),
    .A3(net962),
    .S0(net234),
    .S1(net195),
    .X(net239));
 sky130_fd_sc_hd__and2_1 c324 (.A(net209),
    .B(net239),
    .X(net240));
 sky130_fd_sc_hd__and3_1 c325 (.A(net126),
    .B(net239),
    .C(net729),
    .X(net241));
 sky130_fd_sc_hd__a2111o_1 c326 (.A1(net241),
    .A2(net126),
    .B1(net238),
    .C1(net234),
    .D1(net236),
    .X(net242));
 sky130_fd_sc_hd__buf_1 c327 (.A(net686),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net238),
    .A1(net874),
    .A2(net242),
    .A3(net120),
    .S0(net241),
    .S1(net226),
    .X(net244));
 sky130_fd_sc_hd__and3_1 c329 (.A(net236),
    .B(net232),
    .C(net1061),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c330 (.A(net20),
    .B(net196),
    .C(net114),
    .X(net246));
 sky130_fd_sc_hd__or4bb_1 c331 (.A(net242),
    .B(net92),
    .C_N(net245),
    .D_N(net141),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c332 (.A(net73),
    .B(net958),
    .C(net751),
    .X(net248));
 sky130_fd_sc_hd__and2_1 c333 (.A(net221),
    .B(net685),
    .X(net249));
 sky130_fd_sc_hd__or4bb_1 c334 (.A(net232),
    .B(net246),
    .C_N(net226),
    .D_N(net751),
    .X(net915));
 sky130_fd_sc_hd__sdfrbp_1 c335 (.CLK(clknet_4_9_0_clk),
    .D(net962),
    .RESET_B(net899),
    .SCD(net949),
    .SCE(net751),
    .Q(net251),
    .Q_N(net250));
 sky130_fd_sc_hd__sdfrtn_1 c336 (.CLK_N(clknet_4_9_0_clk),
    .D(net114),
    .RESET_B(net899),
    .SCD(net949),
    .SCE(net998),
    .Q(net252));
 sky130_fd_sc_hd__mux4_2 c337 (.A0(net230),
    .A1(net251),
    .A2(net221),
    .A3(net148),
    .S0(net684),
    .S1(net728),
    .X(net909));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(net873),
    .A1(net141),
    .A2(net243),
    .A3(net144),
    .S0(net879),
    .S1(net949),
    .X(net253));
 sky130_fd_sc_hd__and2_1 c339 (.A(net231),
    .B(net205),
    .X(net254));
 sky130_fd_sc_hd__buf_1 c340 (.A(net737),
    .X(net255));
 sky130_fd_sc_hd__or4bb_1 c341 (.A(net243),
    .B(net234),
    .C_N(net970),
    .D_N(net144),
    .X(net256));
 sky130_fd_sc_hd__sdfrtp_1 c342 (.CLK(clknet_4_2_0_clk),
    .D(net245),
    .RESET_B(net958),
    .SCD(net970),
    .SCE(net242),
    .Q(net257));
 sky130_fd_sc_hd__sdfbbn_1 c343 (.CLK_N(clknet_4_9_0_clk),
    .D(net196),
    .RESET_B(net920),
    .SCD(net230),
    .SCE(net113),
    .SET_B(net970),
    .Q(net259),
    .Q_N(net258));
 sky130_fd_sc_hd__a2111o_1 c344 (.A1(net256),
    .A2(net259),
    .B1(net148),
    .C1(net128),
    .D1(net970),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net256),
    .A1(net257),
    .A2(net970),
    .A3(net949),
    .S0(net250),
    .S1(net966),
    .X(net261));
 sky130_fd_sc_hd__a2111o_2 c346 (.A1(net228),
    .A2(net252),
    .B1(net258),
    .C1(net970),
    .D1(net728),
    .X(net262));
 sky130_fd_sc_hd__sdfbbn_1 c347 (.CLK_N(clknet_4_9_0_clk),
    .D(net257),
    .RESET_B(net909),
    .SCD(net949),
    .SCE(net970),
    .SET_B(net234),
    .Q(net264),
    .Q_N(net263));
 sky130_fd_sc_hd__a2111o_4 c348 (.A1(net264),
    .A2(net221),
    .B1(net258),
    .C1(net825),
    .D1(net734),
    .X(net912));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net260),
    .A1(net949),
    .A2(net254),
    .A3(net234),
    .S0(net912),
    .S1(clknet_1_1__leaf_net752),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net235),
    .A1(net260),
    .A2(net912),
    .A3(net970),
    .S0(net263),
    .S1(net940),
    .X(net266));
 sky130_fd_sc_hd__sdfbbp_1 c351 (.CLK(clknet_4_9_0_clk),
    .D(net970),
    .RESET_B(net912),
    .SCD(net264),
    .SCE(net685),
    .SET_B(net940),
    .Q(net268),
    .Q_N(net267));
 sky130_fd_sc_hd__and3_1 c352 (.A(net228),
    .B(net96),
    .C(net151),
    .X(net269));
 sky130_fd_sc_hd__buf_1 c353 (.A(net726),
    .X(net270));
 sky130_fd_sc_hd__and3_2 c354 (.A(net270),
    .B(net13),
    .C(net148),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 c355 (.A(net726),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 c356 (.A(net724),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net202),
    .A1(net270),
    .A2(net271),
    .A3(net135),
    .S0(net273),
    .S1(net959),
    .X(net274));
 sky130_fd_sc_hd__or4bb_1 c358 (.A(net273),
    .B(net920),
    .C_N(net271),
    .D_N(net734),
    .X(net275));
 sky130_fd_sc_hd__buf_1 c359 (.A(net724),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net272),
    .A1(net937),
    .A2(clknet_1_1__leaf_net154),
    .A3(net968),
    .S0(net872),
    .S1(net940),
    .X(net277));
 sky130_fd_sc_hd__and3_1 c361 (.A(net13),
    .B(net724),
    .C(net940),
    .X(net278));
 sky130_fd_sc_hd__or4bb_4 c362 (.A(net276),
    .B(net96),
    .C_N(net273),
    .D_N(net958),
    .X(net904));
 sky130_fd_sc_hd__and3_1 c363 (.A(net255),
    .B(net276),
    .C(net760),
    .X(net279));
 sky130_fd_sc_hd__or4bb_1 c364 (.A(net958),
    .B(net967),
    .C_N(net35),
    .D_N(clknet_1_1__leaf_net752),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c365 (.A0(net33),
    .A1(net36),
    .A2(net227),
    .A3(net144),
    .S0(clknet_1_0__leaf_net168),
    .S1(net276),
    .X(net281));
 sky130_fd_sc_hd__and3_1 c366 (.A(net251),
    .B(net950),
    .C(net273),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net280),
    .A1(net949),
    .A2(net273),
    .A3(net282),
    .S0(net940),
    .S1(net761),
    .X(net283));
 sky130_fd_sc_hd__sdfbbn_1 c368 (.CLK_N(clknet_4_11_0_clk),
    .D(net269),
    .RESET_B(net36),
    .SCD(clknet_1_0__leaf_net168),
    .SCE(net1060),
    .SET_B(net929),
    .Q(net285),
    .Q_N(net284));
 sky130_fd_sc_hd__and3_1 c369 (.A(net285),
    .B(net927),
    .C(net929),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net148),
    .A1(net927),
    .A2(net92),
    .A3(net925),
    .S0(net269),
    .S1(net940),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net278),
    .A1(net285),
    .A2(net949),
    .A3(net937),
    .S0(net929),
    .S1(net764),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net949),
    .A1(net270),
    .A2(net286),
    .A3(net724),
    .S0(net929),
    .S1(net1058),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net282),
    .A1(net248),
    .A2(net284),
    .A3(net761),
    .S0(net763),
    .S1(net765),
    .X(net290));
 sky130_fd_sc_hd__mux4_2 c392 (.A0(net179),
    .A1(net933),
    .A2(net963),
    .A3(net904),
    .S0(net902),
    .S1(net762),
    .X(net913));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net248),
    .A1(net233),
    .A2(net899),
    .A3(net920),
    .S0(net902),
    .S1(net1055),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net92),
    .A1(net177),
    .A2(net913),
    .A3(net1055),
    .S0(net929),
    .S1(net1047),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net254),
    .A1(net913),
    .A2(net911),
    .S0(net767),
    .S1(net931),
    .X(net293));
 sky130_fd_sc_hd__and2_1 c396 (.A(net972),
    .B(net952),
    .X(net294));
 sky130_fd_sc_hd__dlymetal6s2s_1 c397 (.A(net637),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 c398 (.A(net637),
    .X(net296));
 sky130_fd_sc_hd__and2_1 c399 (.A(net829),
    .B(net71),
    .X(net297));
 sky130_fd_sc_hd__and3_1 c400 (.A(net191),
    .B(net296),
    .C(net195),
    .X(net298));
 sky130_fd_sc_hd__and2_4 c401 (.A(net297),
    .B(net191),
    .X(net886));
 sky130_fd_sc_hd__and2_1 c402 (.A(net297),
    .B(net183),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 c403 (.A(net700),
    .X(net300));
 sky130_fd_sc_hd__buf_1 c404 (.A(net712),
    .X(net301));
 sky130_fd_sc_hd__and2_2 c405 (.A(net301),
    .B(net973),
    .X(net302));
 sky130_fd_sc_hd__and2_1 c406 (.A(net298),
    .B(net195),
    .X(net303));
 sky130_fd_sc_hd__and2_2 c407 (.A(net71),
    .B(net295),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 c408 (.A(net700),
    .X(net916));
 sky130_fd_sc_hd__dlymetal6s2s_1 c409 (.A(net700),
    .X(net305));
 sky130_fd_sc_hd__and2_1 c410 (.A(net305),
    .B(net300),
    .X(net306));
 sky130_fd_sc_hd__mux4_2 c411 (.A0(net306),
    .A1(net295),
    .A2(net305),
    .A3(net301),
    .S0(net297),
    .S1(net973),
    .X(net307));
 sky130_fd_sc_hd__mux4_2 c412 (.A0(net306),
    .A1(net302),
    .A2(net191),
    .A3(net305),
    .S0(net304),
    .S1(net973),
    .X(net308));
 sky130_fd_sc_hd__a2111o_1 c413 (.A1(net305),
    .A2(net303),
    .B1(net306),
    .C1(net304),
    .D1(net973),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net309),
    .A1(net307),
    .A2(net299),
    .A3(net298),
    .S0(net994),
    .S1(net294),
    .X(net310));
 sky130_fd_sc_hd__a2111o_1 c415 (.A1(net298),
    .A2(net305),
    .B1(net836),
    .C1(net307),
    .D1(net309),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 c416 (.A0(net303),
    .A1(net307),
    .A2(net305),
    .A3(net304),
    .S0(net973),
    .S1(net768),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net309),
    .A1(net886),
    .A2(net312),
    .A3(net916),
    .S0(net304),
    .S1(net768),
    .X(net313));
 sky130_fd_sc_hd__and2_0 c418 (.A(net312),
    .B(net220),
    .X(net314));
 sky130_fd_sc_hd__buf_1 c419 (.A(net639),
    .X(net315));
 sky130_fd_sc_hd__and2_0 c420 (.A(net301),
    .B(net899),
    .X(net316));
 sky130_fd_sc_hd__sdfbbn_1 c421 (.CLK_N(clknet_4_0_0_clk),
    .D(net190),
    .RESET_B(net223),
    .SCD(net311),
    .SCE(net839),
    .SET_B(net945),
    .Q(net908),
    .Q_N(net317));
 sky130_fd_sc_hd__a2111o_1 c422 (.A1(net839),
    .A2(net316),
    .B1(net218),
    .C1(net1012),
    .D1(net945),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(net859),
    .A1(net313),
    .A2(net308),
    .A3(net208),
    .S0(net302),
    .S1(net945),
    .X(net319));
 sky130_fd_sc_hd__a2111o_1 c424 (.A1(net220),
    .A2(net86),
    .B1(net302),
    .C1(net945),
    .D1(net223),
    .X(net320));
 sky130_fd_sc_hd__or4bb_1 c425 (.A(net316),
    .B(net89),
    .C_N(net315),
    .D_N(net945),
    .X(net321));
 sky130_fd_sc_hd__sdfrtp_1 c426 (.CLK(clknet_4_0_0_clk),
    .D(net315),
    .RESET_B(net945),
    .SCD(net84),
    .SCE(net711),
    .Q(net322));
 sky130_fd_sc_hd__buf_1 c427 (.A(net638),
    .X(net323));
 sky130_fd_sc_hd__dfbbn_1 c428 (.CLK_N(clknet_4_1_0_clk),
    .D(net218),
    .RESET_B(net946),
    .SET_B(net1041),
    .Q(net325),
    .Q_N(net324));
 sky130_fd_sc_hd__or4bb_1 c429 (.A(net1020),
    .B(net315),
    .C_N(net946),
    .D_N(net738),
    .X(net326));
 sky130_fd_sc_hd__and2_1 c430 (.A(net203),
    .B(net322),
    .X(net327));
 sky130_fd_sc_hd__sdfrtp_1 c431 (.CLK(clknet_4_2_0_clk),
    .D(net944),
    .RESET_B(net1050),
    .SCD(net945),
    .SCE(net740),
    .Q(net328));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net183),
    .A1(net944),
    .A2(net312),
    .A3(net84),
    .S0(net89),
    .S1(net202),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net323),
    .A1(net190),
    .A2(net944),
    .A3(net202),
    .S0(net993),
    .S1(net740),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net323),
    .A1(net944),
    .A2(net312),
    .A3(net697),
    .S0(clknet_1_0__leaf_net769),
    .S1(clknet_1_0__leaf_net770),
    .X(net331));
 sky130_fd_sc_hd__sdfbbp_1 c435 (.CLK(clknet_4_0_0_clk),
    .D(net315),
    .RESET_B(net945),
    .SCD(net301),
    .SCE(net944),
    .SET_B(net996),
    .Q(net333),
    .Q_N(net332));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net333),
    .A1(net205),
    .A2(net916),
    .A3(net944),
    .S0(net1041),
    .S1(clknet_1_1__leaf_net769),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net333),
    .A1(net86),
    .A2(net323),
    .A3(net944),
    .S0(net716),
    .S1(clknet_1_0__leaf_net769),
    .X(net335));
 sky130_fd_sc_hd__buf_2 c438 (.A(net821),
    .X(net336));
 sky130_fd_sc_hd__mux4_2 c439 (.A0(net308),
    .A1(net336),
    .A2(net301),
    .A3(net332),
    .S0(net738),
    .S1(net773),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 c440 (.A(net738),
    .X(net338));
 sky130_fd_sc_hd__and2_0 c441 (.A(net322),
    .B(net120),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 c442 (.A(net738),
    .X(net340));
 sky130_fd_sc_hd__or4bb_1 c443 (.A(net946),
    .B(net866),
    .C_N(net958),
    .D_N(net227),
    .X(net341));
 sky130_fd_sc_hd__and2_0 c444 (.A(net86),
    .B(net129),
    .X(net342));
 sky130_fd_sc_hd__and2_0 c445 (.A(net78),
    .B(net221),
    .X(net343));
 sky130_fd_sc_hd__buf_1 c446 (.A(clknet_1_0__leaf_net744),
    .X(net344));
 sky130_fd_sc_hd__or4bb_1 c447 (.A(net877),
    .B(net78),
    .C_N(net227),
    .D_N(net963),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 c448 (.A(net712),
    .X(net346));
 sky130_fd_sc_hd__sdfbbn_1 c449 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net344),
    .RESET_B(net1045),
    .SCD(net236),
    .SCE(net953),
    .SET_B(net946),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__a2111o_1 c450 (.A1(net236),
    .A2(net835),
    .B1(clknet_1_1__leaf_net344),
    .C1(net954),
    .D1(net302),
    .X(net349));
 sky130_fd_sc_hd__a2111o_4 c451 (.A1(net866),
    .A2(net86),
    .B1(net340),
    .C1(net328),
    .D1(net229),
    .X(net906));
 sky130_fd_sc_hd__or4bb_1 c452 (.A(net345),
    .B(net968),
    .C_N(net322),
    .D_N(clknet_1_1__leaf_net344),
    .X(net350));
 sky130_fd_sc_hd__sdfsbp_1 c453 (.CLK(clknet_4_2_0_clk),
    .D(net1043),
    .SCD(net906),
    .SCE(net205),
    .SET_B(net946),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__a2111o_1 c454 (.A1(net845),
    .A2(net340),
    .B1(clknet_1_1__leaf_net344),
    .C1(net351),
    .D1(net97),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net346),
    .A1(net906),
    .A2(net351),
    .A3(net296),
    .S0(net340),
    .S1(clknet_1_0__leaf_net344),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net873),
    .A1(clknet_1_0__leaf_net353),
    .A2(net97),
    .A3(net906),
    .S0(net345),
    .S1(net240),
    .X(net355));
 sky130_fd_sc_hd__sdfsbp_1 c457 (.CLK(clknet_4_3_0_clk),
    .D(net349),
    .SCD(net352),
    .SCE(clknet_1_1__leaf_net353),
    .SET_B(net774),
    .Q(net357),
    .Q_N(net356));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net835),
    .A1(net352),
    .A2(clknet_1_0__leaf_net350),
    .A3(net946),
    .S0(net774),
    .S1(net776),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 c459 (.A0(clknet_1_0__leaf_net353),
    .A1(net348),
    .A2(net78),
    .A3(net336),
    .S0(clknet_1_0__leaf_net344),
    .S1(net345),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net339),
    .A1(net944),
    .A2(net906),
    .A3(clknet_1_0__leaf_net359),
    .S0(net774),
    .S1(net776),
    .X(net360));
 sky130_fd_sc_hd__a2111o_1 c461 (.A1(clknet_1_0__leaf_net359),
    .A2(net239),
    .B1(net347),
    .C1(net845),
    .X(net361));
 sky130_fd_sc_hd__and2_0 c462 (.A(net268),
    .B(net302),
    .X(net362));
 sky130_fd_sc_hd__and2_1 c463 (.A(net302),
    .B(net899),
    .X(net363));
 sky130_fd_sc_hd__and2_0 c464 (.A(net252),
    .B(net886),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 c465 (.A(net635),
    .X(net365));
 sky130_fd_sc_hd__and2_0 c466 (.A(net246),
    .B(net268),
    .X(net366));
 sky130_fd_sc_hd__and2_0 c467 (.A(net365),
    .B(net135),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net635),
    .X(net368));
 sky130_fd_sc_hd__and2_0 c469 (.A(net113),
    .B(net268),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net912),
    .A1(net317),
    .A2(net195),
    .A3(net363),
    .S0(net956),
    .S1(net737),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net141),
    .A1(net841),
    .A2(net906),
    .A3(net975),
    .S0(net956),
    .S1(net901),
    .X(net371));
 sky130_fd_sc_hd__and2_0 c472 (.A(clknet_1_0__leaf_net350),
    .B(net901),
    .X(net372));
 sky130_fd_sc_hd__and2_0 c473 (.A(net367),
    .B(clknet_1_0__leaf_net372),
    .X(net373));
 sky130_fd_sc_hd__a2111o_1 c474 (.A1(net366),
    .A2(net883),
    .B1(net252),
    .C1(net190),
    .D1(net956),
    .X(net374));
 sky130_fd_sc_hd__or4bb_1 c475 (.A(net234),
    .B(net867),
    .C_N(net956),
    .D_N(net901),
    .X(net375));
 sky130_fd_sc_hd__and2_0 c476 (.A(clknet_1_0__leaf_net373),
    .B(net901),
    .X(net376));
 sky130_fd_sc_hd__sdfstp_1 c477 (.CLK(clknet_4_9_0_clk),
    .D(net375),
    .SCD(clknet_1_0__leaf_net376),
    .SCE(net956),
    .SET_B(net1039),
    .Q(net377));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net369),
    .A1(net240),
    .A2(net956),
    .A3(clknet_1_1__leaf_net350),
    .S0(net267),
    .S1(clknet_1_1__leaf_net373),
    .X(net378));
 sky130_fd_sc_hd__and3_2 c479 (.A(net226),
    .B(net375),
    .C(net956),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net195),
    .A1(net363),
    .A2(net375),
    .A3(net336),
    .S0(net141),
    .S1(net377),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net227),
    .A1(net313),
    .A2(net956),
    .A3(net351),
    .S0(net775),
    .S1(net779),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net376),
    .A1(net895),
    .A2(net356),
    .A3(net363),
    .S0(clknet_1_0__leaf_net373),
    .S1(net779),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net378),
    .A1(net834),
    .A2(clknet_1_1__leaf_net350),
    .A3(net336),
    .S0(net363),
    .S1(net267),
    .X(net382));
 sky130_fd_sc_hd__a2111o_1 c484 (.A1(net262),
    .A2(clknet_1_0__leaf_net887),
    .B1(net895),
    .C1(clknet_1_0__leaf_net168),
    .D1(net958),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(clknet_1_1__leaf_net168),
    .A1(net956),
    .A2(net202),
    .A3(net950),
    .S0(net716),
    .S1(net761),
    .X(net384));
 sky130_fd_sc_hd__sdfbbn_1 c486 (.CLK_N(clknet_4_14_0_clk),
    .D(net959),
    .RESET_B(net286),
    .SCD(net920),
    .SCE(net135),
    .SET_B(net767),
    .Q(net386),
    .Q_N(net385));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net279),
    .A1(clknet_1_1__leaf_net168),
    .A2(net385),
    .A3(net262),
    .S0(net967),
    .S1(net765),
    .X(net387));
 sky130_fd_sc_hd__sdfbbp_1 c488 (.CLK(clknet_4_11_0_clk),
    .D(net13),
    .RESET_B(net271),
    .SCD(net286),
    .SCE(net901),
    .SET_B(net1036),
    .Q(net389),
    .Q_N(net388));
 sky130_fd_sc_hd__a2111o_1 c489 (.A1(net904),
    .A2(net279),
    .B1(net223),
    .C1(net761),
    .D1(net1033),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net273),
    .A1(net388),
    .A2(clknet_1_1__leaf_net887),
    .A3(net271),
    .S0(net227),
    .S1(net950),
    .X(net391));
 sky130_fd_sc_hd__sdfbbn_1 c491 (.CLK_N(clknet_4_9_0_clk),
    .D(net970),
    .RESET_B(net848),
    .SCD(net912),
    .SCE(net920),
    .SET_B(net952),
    .Q(net393),
    .Q_N(net392));
 sky130_fd_sc_hd__a2111o_1 c492 (.A1(net389),
    .A2(net392),
    .B1(net958),
    .C1(clknet_1_1__leaf_net887),
    .D1(net766),
    .X(net919));
 sky130_fd_sc_hd__mux4_2 c493 (.A0(net286),
    .A1(net389),
    .A2(net336),
    .A3(net954),
    .S0(net968),
    .S1(net780),
    .X(net394));
 sky130_fd_sc_hd__sdfbbn_1 c494 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net168),
    .RESET_B(net394),
    .SCD(clknet_1_0__leaf_net919),
    .SCE(net904),
    .SET_B(net781),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__a2111o_1 c495 (.A1(net394),
    .A2(net273),
    .B1(net916),
    .C1(net690),
    .D1(net1036),
    .X(net397));
 sky130_fd_sc_hd__a2111o_1 c496 (.A1(net374),
    .A2(net392),
    .B1(net1063),
    .C1(net959),
    .D1(net1032),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net872),
    .A1(net135),
    .A2(net984),
    .A3(net886),
    .S0(net968),
    .S1(net719),
    .X(net399));
 sky130_fd_sc_hd__a2111o_2 c498 (.A1(net399),
    .A2(net395),
    .B1(net273),
    .C1(net696),
    .D1(net726),
    .X(net400));
 sky130_fd_sc_hd__a2111o_1 c499 (.A1(net225),
    .A2(net394),
    .B1(net1057),
    .C1(net286),
    .D1(net967),
    .X(net401));
 sky130_fd_sc_hd__a2111o_1 c500 (.A1(net161),
    .A2(net959),
    .B1(net279),
    .C1(net286),
    .D1(net1053),
    .X(net402));
 sky130_fd_sc_hd__sdfbbp_1 c501 (.CLK(clknet_4_14_0_clk),
    .D(net249),
    .RESET_B(net402),
    .SCD(net920),
    .SCE(net394),
    .SET_B(net1037),
    .Q(net404),
    .Q_N(net403));
 sky130_fd_sc_hd__a2111o_1 c502 (.A1(net396),
    .A2(net336),
    .B1(net394),
    .C1(net1009),
    .D1(net780),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net227),
    .A1(net279),
    .A2(net144),
    .A3(net886),
    .S0(net403),
    .S1(net917),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net352),
    .A1(net336),
    .A2(net404),
    .A3(net395),
    .S0(net920),
    .S1(net734),
    .X(net407));
 sky130_fd_sc_hd__a2111o_1 c505 (.A1(net406),
    .A2(net867),
    .B1(clknet_1_0__leaf_net919),
    .C1(net29),
    .D1(net403),
    .X(net889));
 sky130_fd_sc_hd__and2_1 c528 (.A(net299),
    .B(net834),
    .X(net408));
 sky130_fd_sc_hd__buf_2 c529 (.A(net1028),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 c530 (.A(net702),
    .X(net410));
 sky130_fd_sc_hd__and2_2 c531 (.A(net307),
    .B(net409),
    .X(net411));
 sky130_fd_sc_hd__and2_1 c532 (.A(net411),
    .B(net300),
    .X(net412));
 sky130_fd_sc_hd__and2_0 c533 (.A(net974),
    .B(net299),
    .X(net413));
 sky130_fd_sc_hd__and2_1 c534 (.A(net413),
    .B(net412),
    .X(net414));
 sky130_fd_sc_hd__and2_1 c535 (.A(net413),
    .B(net409),
    .X(net415));
 sky130_fd_sc_hd__and2_0 c536 (.A(net414),
    .B(net412),
    .X(net416));
 sky130_fd_sc_hd__and2_0 c537 (.A(net68),
    .B(net410),
    .X(net417));
 sky130_fd_sc_hd__a2111o_2 c538 (.A1(net408),
    .A2(net886),
    .B1(net413),
    .C1(net411),
    .D1(net414),
    .X(net418));
 sky130_fd_sc_hd__or4bb_1 c539 (.A(net300),
    .B(net295),
    .C_N(net411),
    .D_N(net409),
    .X(net419));
 sky130_fd_sc_hd__and2_0 c540 (.A(net835),
    .B(net916),
    .X(net420));
 sky130_fd_sc_hd__and2_0 c541 (.A(net416),
    .B(net414),
    .X(net421));
 sky130_fd_sc_hd__and2_0 c542 (.A(net414),
    .B(net415),
    .X(net422));
 sky130_fd_sc_hd__a2111o_1 c543 (.A1(net419),
    .A2(net952),
    .B1(net1008),
    .C1(net414),
    .D1(net422),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(net410),
    .A1(net421),
    .A2(net412),
    .A3(net423),
    .S0(net409),
    .S1(net974),
    .X(net424));
 sky130_fd_sc_hd__or4bb_1 c545 (.A(net422),
    .B(net420),
    .C_N(net997),
    .D_N(net784),
    .X(net425));
 sky130_fd_sc_hd__or4bb_1 c546 (.A(net916),
    .B(net423),
    .C_N(net425),
    .D_N(net785),
    .X(net426));
 sky130_fd_sc_hd__a2111o_1 c547 (.A1(net423),
    .A2(net72),
    .B1(net411),
    .D1(net784),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c548 (.A0(net425),
    .A1(net419),
    .A2(net417),
    .A3(net423),
    .S0(net952),
    .S1(net414),
    .X(net428));
 sky130_fd_sc_hd__or4bb_2 c549 (.A(net624),
    .B(net75),
    .C_N(net679),
    .D_N(net786),
    .X(net429));
 sky130_fd_sc_hd__buf_1 c550 (.A(net641),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(net206),
    .A1(net324),
    .A2(net418),
    .A3(net205),
    .S0(net946),
    .S1(net768),
    .X(net431));
 sky130_fd_sc_hd__and2_0 c552 (.A(net325),
    .B(net768),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c553 (.A(net641),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 c554 (.A(net739),
    .X(net434));
 sky130_fd_sc_hd__buf_1 c555 (.A(net739),
    .X(net435));
 sky130_fd_sc_hd__and3_1 c556 (.A(net433),
    .B(net218),
    .C(net689),
    .X(net436));
 sky130_fd_sc_hd__and2_0 c557 (.A(net961),
    .B(net768),
    .X(net437));
 sky130_fd_sc_hd__and2_0 c558 (.A(net409),
    .B(net689),
    .X(net438));
 sky130_fd_sc_hd__or4bb_2 c559 (.A(net436),
    .B(net218),
    .C_N(net961),
    .D_N(net969),
    .X(net893));
 sky130_fd_sc_hd__or4bb_1 c560 (.A(net218),
    .B(net960),
    .C_N(net437),
    .D_N(net945),
    .X(net439));
 sky130_fd_sc_hd__and2_0 c561 (.A(net434),
    .B(net960),
    .X(net440));
 sky130_fd_sc_hd__or4bb_4 c562 (.A(net408),
    .B(net205),
    .C_N(net961),
    .D_N(net960),
    .X(net441));
 sky130_fd_sc_hd__or4bb_1 c563 (.A(net432),
    .B(net969),
    .C_N(net437),
    .D_N(clknet_1_0__leaf_net771),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 c564 (.A(net739),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c565 (.A(net443),
    .B(net886),
    .C(net441),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net442),
    .A1(net441),
    .A2(net438),
    .A3(net430),
    .S0(net444),
    .S1(net433),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c567 (.A(clknet_1_1__leaf_net445),
    .B(net444),
    .C(net440),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(clknet_1_0__leaf_net446),
    .A1(net408),
    .A2(net441),
    .A3(clknet_1_0__leaf_net445),
    .S0(net969),
    .S1(net960),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 c569 (.A(net820),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net420),
    .A1(net448),
    .A2(net443),
    .A3(net960),
    .S0(clknet_1_1__leaf_net446),
    .S1(net787),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net437),
    .A1(clknet_1_0__leaf_net446),
    .A2(net444),
    .A3(net969),
    .S0(net787),
    .S1(net971),
    .X(net450));
 sky130_fd_sc_hd__sdfbbn_1 c572 (.CLK_N(clknet_4_3_0_clk),
    .D(net448),
    .RESET_B(clknet_1_1__leaf_net359),
    .SCD(net347),
    .SCE(net705),
    .SET_B(net758),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__a2111o_1 c573 (.A1(net409),
    .A2(net452),
    .B1(clknet_1_1__leaf_net359),
    .C1(net961),
    .D1(net948),
    .X(net453));
 sky130_fd_sc_hd__or4bb_2 c574 (.A(net452),
    .B(net871),
    .C_N(net953),
    .D_N(net775),
    .X(net454));
 sky130_fd_sc_hd__or4bb_1 c575 (.A(net1031),
    .B(net947),
    .C_N(net451),
    .D_N(net202),
    .X(net455));
 sky130_fd_sc_hd__or4bb_1 c576 (.A(net229),
    .B(net871),
    .C_N(net969),
    .D_N(net960),
    .X(net456));
 sky130_fd_sc_hd__sdfbbn_1 c577 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net359),
    .RESET_B(net68),
    .SCD(net874),
    .SCE(net229),
    .SET_B(net429),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__or4bb_1 c578 (.A(net342),
    .B(net409),
    .C_N(net963),
    .D_N(net777),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 c579 (.A0(net239),
    .A1(net960),
    .A2(net863),
    .A3(net348),
    .S0(net836),
    .S1(net886),
    .X(net460));
 sky130_fd_sc_hd__a2111o_1 c580 (.A1(net237),
    .A2(net458),
    .B1(net454),
    .C1(net955),
    .D1(net683),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net448),
    .A1(net457),
    .A2(net948),
    .A3(net689),
    .S0(clknet_1_0__leaf_net707),
    .S1(net774),
    .X(net462));
 sky130_fd_sc_hd__a2111o_1 c582 (.A1(net863),
    .A2(net874),
    .B1(net458),
    .C1(net1031),
    .D1(net953),
    .X(net463));
 sky130_fd_sc_hd__a2111o_1 c583 (.A1(net208),
    .A2(net961),
    .B1(net960),
    .C1(net971),
    .D1(clknet_1_0__leaf_net884),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net836),
    .A1(net452),
    .A2(net68),
    .A3(net448),
    .S0(net948),
    .S1(clknet_1_0__leaf_net884),
    .X(net465));
 sky130_fd_sc_hd__sdfbbp_1 c585 (.CLK(clknet_4_3_0_clk),
    .D(net1046),
    .RESET_B(net463),
    .SCD(net296),
    .SCE(net704),
    .SET_B(clknet_1_0__leaf_net884),
    .Q(net467),
    .Q_N(net466));
 sky130_fd_sc_hd__a2111o_1 c586 (.A1(clknet_1_1__leaf_net464),
    .A2(net458),
    .B1(net125),
    .C1(net706),
    .D1(clknet_1_0__leaf_net884),
    .X(net468));
 sky130_fd_sc_hd__a2111o_1 c587 (.A1(net296),
    .A2(clknet_1_0__leaf_net464),
    .B1(net955),
    .C1(net467),
    .D1(clknet_1_0__leaf_net884),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net348),
    .A1(net468),
    .A2(clknet_1_0__leaf_net464),
    .A3(net451),
    .S0(net961),
    .S1(net466),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 c589 (.A0(net415),
    .A1(net467),
    .A2(net89),
    .A3(net229),
    .S0(net463),
    .S1(net451),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net463),
    .A1(clknet_1_0__leaf_net464),
    .A2(clknet_1_0__leaf_net359),
    .A3(net454),
    .S0(net955),
    .S1(net759),
    .X(net472));
 sky130_fd_sc_hd__sdfbbn_1 c591 (.CLK_N(clknet_4_3_0_clk),
    .D(net459),
    .RESET_B(net456),
    .SCD(net463),
    .SCE(net961),
    .SET_B(net867),
    .Q(net474),
    .Q_N(net473));
 sky130_fd_sc_hd__sdfbbn_1 c592 (.CLK_N(clknet_4_3_0_clk),
    .D(net1042),
    .RESET_B(net441),
    .SCD(clknet_1_1__leaf_net464),
    .SCE(clknet_1_0__leaf_net469),
    .SET_B(net1048),
    .Q(net476),
    .Q_N(net475));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net237),
    .A1(clknet_1_1__leaf_net464),
    .A2(net476),
    .A3(net457),
    .S0(net473),
    .S1(net706),
    .X(net477));
 sky130_fd_sc_hd__and3_1 c594 (.A(net129),
    .B(net893),
    .C(net706),
    .X(net478));
 sky130_fd_sc_hd__and3_1 c595 (.A(net362),
    .B(net129),
    .C(net457),
    .X(net479));
 sky130_fd_sc_hd__or4bb_1 c596 (.A(net205),
    .B(net135),
    .C_N(net957),
    .D_N(clknet_1_0__leaf_net884),
    .X(net480));
 sky130_fd_sc_hd__and3_1 c597 (.A(net479),
    .B(net259),
    .C(net834),
    .X(net481));
 sky130_fd_sc_hd__and3_1 c598 (.A(clknet_1_1__leaf_net480),
    .B(net957),
    .C(net258),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 c599 (.A(net818),
    .X(net483));
 sky130_fd_sc_hd__a2111o_1 c600 (.A1(net377),
    .A2(clknet_1_0__leaf_net480),
    .B1(net479),
    .C1(net435),
    .D1(net957),
    .X(net484));
 sky130_fd_sc_hd__or4bb_2 c601 (.A(net483),
    .B(net867),
    .C_N(net13),
    .D_N(net135),
    .X(net485));
 sky130_fd_sc_hd__a2111o_1 c602 (.A1(net961),
    .A2(net953),
    .B1(net13),
    .C1(net485),
    .D1(net969),
    .X(net486));
 sky130_fd_sc_hd__sdfbbp_1 c603 (.CLK(clknet_4_3_0_clk),
    .D(net486),
    .RESET_B(net476),
    .SCD(clknet_1_0__leaf_net480),
    .SCE(net775),
    .SET_B(clknet_1_0__leaf_net789),
    .Q(net942),
    .Q_N(net487));
 sky130_fd_sc_hd__a2111o_1 c604 (.A1(net942),
    .A2(net475),
    .B1(net963),
    .C1(net961),
    .D1(net706),
    .X(net488));
 sky130_fd_sc_hd__sdfstp_1 c605 (.CLK(clknet_4_12_0_clk),
    .D(net488),
    .SCD(net486),
    .SCE(net475),
    .SET_B(net895),
    .Q(net489));
 sky130_fd_sc_hd__and3_1 c606 (.A(net953),
    .B(net135),
    .C(net1030),
    .X(net490));
 sky130_fd_sc_hd__a2111o_1 c607 (.A1(net490),
    .A2(net1030),
    .B1(net1035),
    .C1(net1065),
    .D1(net481),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net485),
    .A1(net486),
    .A2(net488),
    .A3(net674),
    .S0(net682),
    .S1(clknet_1_0__leaf_net770),
    .X(net492));
 sky130_fd_sc_hd__a2111o_1 c609 (.A1(net430),
    .A2(net942),
    .B1(net673),
    .C1(clknet_1_1__leaf_net884),
    .D1(clknet_1_0__leaf_net892),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net125),
    .A1(net488),
    .A2(net240),
    .A3(net221),
    .S0(net481),
    .S1(net955),
    .X(net493));
 sky130_fd_sc_hd__a2111o_1 c611 (.A1(net259),
    .A2(clknet_1_1__leaf_net469),
    .B1(net871),
    .C1(net775),
    .D1(net778),
    .X(net494));
 sky130_fd_sc_hd__sdfbbn_1 c612 (.CLK_N(clknet_4_6_0_clk),
    .D(net493),
    .RESET_B(net488),
    .SCD(net486),
    .SCE(net490),
    .SET_B(net485),
    .Q(net496),
    .Q_N(net495));
 sky130_fd_sc_hd__or4bb_2 c613 (.A(net476),
    .B(net495),
    .C_N(net377),
    .D_N(net674),
    .X(net497));
 sky130_fd_sc_hd__and3_1 c614 (.A(net496),
    .B(net1030),
    .C(net689),
    .X(net498));
 sky130_fd_sc_hd__sdfbbn_1 c615 (.CLK_N(clknet_4_6_0_clk),
    .D(net240),
    .RESET_B(net498),
    .SCD(net489),
    .SCE(net486),
    .SET_B(clknet_1_0__leaf_net892),
    .Q(net500),
    .Q_N(net499));
 sky130_fd_sc_hd__mux4_2 c616 (.A0(net969),
    .A1(net400),
    .A2(net404),
    .A3(net386),
    .S0(net777),
    .S1(net778),
    .X(net501));
 sky130_fd_sc_hd__mux4_2 c617 (.A0(net485),
    .A1(net400),
    .A2(net457),
    .A3(net767),
    .S0(net776),
    .S1(net782),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net151),
    .A1(net393),
    .A2(net502),
    .A3(net848),
    .S0(net950),
    .S1(net998),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net953),
    .A1(net957),
    .A2(net950),
    .A3(net848),
    .S0(net777),
    .S1(clknet_1_1__leaf_net789),
    .X(net504));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net840),
    .A1(net842),
    .A2(net3),
    .A3(net866),
    .S0(net875),
    .S1(net868),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net404),
    .A1(net357),
    .A2(clknet_1_0__leaf_net889),
    .A3(net969),
    .S0(net916),
    .S1(net938),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net271),
    .A1(net31),
    .A2(net144),
    .A3(net927),
    .S0(net957),
    .S1(clknet_1_0__leaf_net889),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net489),
    .A1(net1007),
    .A2(net886),
    .A3(net404),
    .S0(net953),
    .S1(clknet_1_1__leaf_net770),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net89),
    .A1(net1009),
    .A2(net916),
    .A3(net502),
    .S0(net927),
    .S1(clknet_1_0__leaf_net887),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net368),
    .A1(net501),
    .A2(net893),
    .A3(net403),
    .S0(net233),
    .S1(net777),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net393),
    .A1(net927),
    .A2(net123),
    .A3(net31),
    .S0(net954),
    .S1(net780),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net458),
    .A1(net963),
    .A2(net969),
    .A3(clknet_1_0__leaf_net507),
    .S0(clknet_1_1__leaf_net770),
    .S1(clknet_1_0__leaf_net892),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net504),
    .A1(net271),
    .A2(net927),
    .A3(net487),
    .S0(clknet_1_0__leaf_net887),
    .S1(net791),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net957),
    .A1(clknet_1_1__leaf_net507),
    .A2(net938),
    .A3(net13),
    .S0(net135),
    .S1(net767),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net510),
    .A1(net202),
    .A2(net400),
    .A3(net271),
    .S0(net778),
    .S1(net794),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net877),
    .A1(net840),
    .A2(net875),
    .A3(net0),
    .S0(net861),
    .S1(net828),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net386),
    .A1(net123),
    .A2(net403),
    .A3(clknet_1_0__leaf_net710),
    .S0(net767),
    .S1(net794),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net135),
    .A1(net502),
    .A2(net123),
    .A3(net780),
    .S0(clknet_1_0__leaf_net892),
    .S1(net897),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_0__leaf_net507),
    .A1(net400),
    .A2(net703),
    .A3(net792),
    .S0(net794),
    .S1(net795),
    .X(net517));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net357),
    .A1(net404),
    .A2(net502),
    .A3(net886),
    .S0(net790),
    .S1(net794),
    .X(net518));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_1__leaf_net507),
    .A1(net832),
    .A2(net969),
    .A3(clknet_1_0__leaf_net887),
    .S0(net694),
    .S1(net795),
    .X(net519));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net144),
    .A1(net938),
    .A2(net788),
    .A3(net793),
    .S0(net794),
    .S1(net797),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net515),
    .A1(net938),
    .A2(clknet_1_1__leaf_net710),
    .A3(clknet_1_1__leaf_net884),
    .S0(net794),
    .S1(net797),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net867),
    .A1(net520),
    .A2(net501),
    .A3(net734),
    .S0(net767),
    .S1(net1054),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net863),
    .A1(net842),
    .A2(net864),
    .A3(net870),
    .S0(net0),
    .S1(net845),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net878),
    .A1(net848),
    .A2(net851),
    .A3(net825),
    .S0(net836),
    .S1(net841),
    .X(net3));
 sky130_fd_sc_hd__and2_0 c66 (.A(net825),
    .B(net830),
    .X(net4));
 sky130_fd_sc_hd__and2_1 c660 (.A(net67),
    .B(net304),
    .X(net523));
 sky130_fd_sc_hd__and2_1 c661 (.A(net304),
    .B(net412),
    .X(net524));
 sky130_fd_sc_hd__and2_2 c662 (.A(net412),
    .B(net784),
    .X(net525));
 sky130_fd_sc_hd__and2_2 c663 (.A(net304),
    .B(net525),
    .X(net526));
 sky130_fd_sc_hd__and2_4 c664 (.A(net525),
    .B(net524),
    .X(net527));
 sky130_fd_sc_hd__and2_1 c665 (.A(net416),
    .B(net834),
    .X(net528));
 sky130_fd_sc_hd__and2_1 c666 (.A(net768),
    .B(net786),
    .X(net529));
 sky130_fd_sc_hd__and2_2 c667 (.A(net85),
    .B(net524),
    .X(net530));
 sky130_fd_sc_hd__and2_1 c668 (.A(net525),
    .B(net529),
    .X(net531));
 sky130_fd_sc_hd__or4bb_1 c669 (.A(net525),
    .B(net529),
    .C_N(net785),
    .D_N(net786),
    .X(net532));
 sky130_fd_sc_hd__and2_1 c67 (.A(net841),
    .B(net834),
    .X(net5));
 sky130_fd_sc_hd__and2_1 c670 (.A(net72),
    .B(net531),
    .X(net533));
 sky130_fd_sc_hd__and2_0 c671 (.A(net307),
    .B(net525),
    .X(net534));
 sky130_fd_sc_hd__and2_0 c672 (.A(net534),
    .B(net533),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net530),
    .A1(net527),
    .A2(net525),
    .A3(net528),
    .S0(net411),
    .S1(net785),
    .X(net536));
 sky130_fd_sc_hd__and3_1 c674 (.A(net421),
    .B(net412),
    .C(net530),
    .X(net537));
 sky130_fd_sc_hd__and3_1 c675 (.A(net536),
    .B(net988),
    .C(net786),
    .X(net538));
 sky130_fd_sc_hd__and3_1 c676 (.A(net536),
    .B(net530),
    .C(net537),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 c677 (.A(net1028),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net535),
    .A1(net528),
    .A2(net536),
    .A3(net538),
    .S0(net527),
    .S1(net537),
    .X(net541));
 sky130_fd_sc_hd__buf_1 c679 (.A(net1028),
    .X(net542));
 sky130_fd_sc_hd__and2_1 c68 (.A(net865),
    .B(net871),
    .X(net6));
 sky130_fd_sc_hd__and3_1 c680 (.A(net533),
    .B(net536),
    .C(net418),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net540),
    .A1(net543),
    .A2(net542),
    .A3(net536),
    .S0(net525),
    .S1(net532),
    .X(net544));
 sky130_fd_sc_hd__sdfstp_2 c682 (.CLK(clknet_4_5_0_clk),
    .D(net542),
    .SCD(net441),
    .SCE(net947),
    .SET_B(net1034),
    .Q(net545));
 sky130_fd_sc_hd__and3_1 c683 (.A(net85),
    .B(net532),
    .C(net222),
    .X(net546));
 sky130_fd_sc_hd__or4bb_1 c684 (.A(net222),
    .B(net527),
    .C_N(net530),
    .D_N(net732),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 c685 (.A(net740),
    .X(net548));
 sky130_fd_sc_hd__and3_1 c686 (.A(net444),
    .B(net411),
    .C(net732),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net539),
    .A1(net547),
    .A2(net528),
    .A3(net545),
    .S0(net947),
    .S1(net1044),
    .X(net550));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net337),
    .A1(net1010),
    .A2(net222),
    .A3(net947),
    .S0(net539),
    .S1(net542),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 c689 (.A(net740),
    .X(net552));
 sky130_fd_sc_hd__and2_1 c69 (.A(net2),
    .B(net6),
    .X(net7));
 sky130_fd_sc_hd__sdfbbp_1 c690 (.CLK(clknet_4_4_0_clk),
    .D(net548),
    .RESET_B(net543),
    .SCD(net545),
    .SCE(net441),
    .SET_B(net947),
    .Q(net554),
    .Q_N(net553));
 sky130_fd_sc_hd__or4bb_2 c691 (.A(net553),
    .B(net444),
    .C_N(net680),
    .D_N(net787),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net85),
    .A1(net444),
    .A2(net528),
    .A3(net548),
    .S0(net555),
    .S1(net699),
    .X(net556));
 sky130_fd_sc_hd__sedfxbp_1 c693 (.CLK(clknet_4_5_0_clk),
    .D(net549),
    .DE(net991),
    .SCD(net542),
    .SCE(net947),
    .Q(net558),
    .Q_N(net557));
 sky130_fd_sc_hd__and3_2 c694 (.A(net552),
    .B(net768),
    .C(net800),
    .X(net559));
 sky130_fd_sc_hd__and3_1 c695 (.A(net558),
    .B(net526),
    .C(net559),
    .X(net560));
 sky130_fd_sc_hd__or4bb_4 c696 (.A(net532),
    .B(net337),
    .C_N(net557),
    .D_N(net787),
    .X(net561));
 sky130_fd_sc_hd__or4bb_2 c697 (.A(net528),
    .B(net559),
    .C_N(net951),
    .D_N(net531),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net537),
    .A1(net85),
    .A2(net562),
    .A3(net559),
    .S0(net951),
    .S1(net971),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(net418),
    .A1(net954),
    .A2(net562),
    .A3(net559),
    .S0(net971),
    .S1(net1056),
    .X(net564));
 sky130_fd_sc_hd__and3_1 c70 (.A(net864),
    .B(net871),
    .C(net825),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net560),
    .A1(net559),
    .A2(net562),
    .A3(net699),
    .S0(net802),
    .S1(net803),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net547),
    .A1(net555),
    .A2(net526),
    .A3(net529),
    .S0(net562),
    .S1(clknet_1_1__leaf_net744),
    .X(net566));
 sky130_fd_sc_hd__mux4_2 c702 (.A0(net523),
    .A1(net418),
    .A2(net951),
    .A3(net559),
    .S0(clknet_1_1__leaf_net744),
    .S1(net803),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net562),
    .A1(net545),
    .A2(clknet_1_0__leaf_net567),
    .A3(net555),
    .S0(net527),
    .S1(net699),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 c704 (.A(net815),
    .X(net569));
 sky130_fd_sc_hd__or4bb_4 c705 (.A(clknet_1_0__leaf_net567),
    .B(net545),
    .C_N(net441),
    .D_N(net556),
    .X(net570));
 sky130_fd_sc_hd__a2111o_1 c706 (.A1(net569),
    .A2(clknet_1_0__leaf_net477),
    .B1(net223),
    .C1(net948),
    .D1(net971),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net815),
    .X(net572));
 sky130_fd_sc_hd__and3_1 c708 (.A(net572),
    .B(net883),
    .C(net971),
    .X(net573));
 sky130_fd_sc_hd__and3_1 c709 (.A(net554),
    .B(clknet_1_0__leaf_net708),
    .C(net971),
    .X(net574));
 sky130_fd_sc_hd__and2_1 c71 (.A(net8),
    .B(net872),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 c710 (.A(net739),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net555),
    .A1(net575),
    .A2(net951),
    .A3(net868),
    .S0(net120),
    .S1(net955),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 c712 (.A(net821),
    .X(net577));
 sky130_fd_sc_hd__sdfbbn_1 c713 (.CLK_N(clknet_4_5_0_clk),
    .D(net529),
    .RESET_B(clknet_1_1__leaf_net477),
    .SCD(net947),
    .SCE(net962),
    .SET_B(net411),
    .Q(net579),
    .Q_N(net578));
 sky130_fd_sc_hd__buf_1 c714 (.A(clknet_1_0__leaf_net744),
    .X(net580));
 sky130_fd_sc_hd__sedfxbp_1 c715 (.CLK(clknet_4_5_0_clk),
    .D(net576),
    .DE(net531),
    .SCD(net523),
    .SCE(net952),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__and3_1 c716 (.A(net411),
    .B(net575),
    .C(net581),
    .X(net583));
 sky130_fd_sc_hd__a2111o_2 c717 (.A1(net120),
    .A2(net530),
    .B1(net441),
    .C1(net997),
    .D1(net559),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net559),
    .A1(net580),
    .A2(net989),
    .A3(net583),
    .S0(net101),
    .S1(net584),
    .X(net585));
 sky130_fd_sc_hd__and3_1 c719 (.A(net531),
    .B(net951),
    .C(net962),
    .X(net586));
 sky130_fd_sc_hd__and3_1 c72 (.A(net871),
    .B(net1),
    .C(net2),
    .X(net10));
 sky130_fd_sc_hd__and3_1 c720 (.A(net573),
    .B(net584),
    .C(net578),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net538),
    .A1(net411),
    .A2(net583),
    .A3(net584),
    .S0(net340),
    .S1(net530),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net523),
    .A1(net582),
    .A2(net586),
    .A3(clknet_1_1__leaf_net567),
    .S0(net955),
    .S1(net951),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net586),
    .A1(net584),
    .A2(net454),
    .A3(net803),
    .S0(net805),
    .S1(clknet_1_0__leaf_net806),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net546),
    .A1(net586),
    .A2(net947),
    .A3(net543),
    .S0(net717),
    .S1(clknet_1_0__leaf_net806),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 c725 (.A(net1052),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net868),
    .A1(net951),
    .A2(net989),
    .A3(net733),
    .S0(net788),
    .S1(clknet_1_0__leaf_net806),
    .X(net593));
 sky130_fd_sc_hd__sedfxtp_4 c727 (.CLK(clknet_4_6_0_clk),
    .D(net221),
    .DE(net593),
    .SCD(net581),
    .SCE(net13),
    .Q(net594));
 sky130_fd_sc_hd__a2111o_1 c728 (.A1(net834),
    .A2(net340),
    .B1(clknet_1_1__leaf_net372),
    .C1(net584),
    .D1(net805),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net951),
    .A1(net579),
    .A2(net526),
    .A3(net340),
    .S0(net955),
    .S1(net804),
    .X(net596));
 sky130_fd_sc_hd__and2_1 c73 (.A(net10),
    .B(net8),
    .X(net11));
 sky130_fd_sc_hd__or4bb_1 c730 (.A(net584),
    .B(net596),
    .C_N(net867),
    .D_N(net594),
    .X(net597));
 sky130_fd_sc_hd__a2111o_1 c731 (.A1(net484),
    .A2(net545),
    .B1(net963),
    .C1(net594),
    .D1(net575),
    .X(net598));
 sky130_fd_sc_hd__a2111o_1 c732 (.A1(net951),
    .A2(net584),
    .B1(net594),
    .C1(net441),
    .D1(net955),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net441),
    .A1(net582),
    .A2(net943),
    .A3(net594),
    .S0(net867),
    .S1(net805),
    .X(net600));
 sky130_fd_sc_hd__sdfbbn_1 c734 (.CLK_N(clknet_4_7_0_clk),
    .D(net583),
    .RESET_B(net594),
    .SCD(net527),
    .SCE(net340),
    .SET_B(net943),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__sdfbbp_1 c735 (.CLK(clknet_4_7_0_clk),
    .D(net340),
    .RESET_B(net592),
    .SCD(net943),
    .SCE(clknet_1_0__leaf_net595),
    .SET_B(net601),
    .Q(net603));
 sky130_fd_sc_hd__a2111o_1 c736 (.A1(net955),
    .A2(net602),
    .B1(net943),
    .C1(net340),
    .D1(net1059),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_0__leaf_net372),
    .A1(net497),
    .A2(net599),
    .A3(net578),
    .S0(net955),
    .S1(net799),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net990),
    .A1(net594),
    .A2(net601),
    .A3(net599),
    .S0(net714),
    .S1(net735),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net478),
    .A1(net602),
    .A2(net460),
    .A3(net943),
    .S0(net497),
    .S1(net805),
    .X(net607));
 sky130_fd_sc_hd__and2_0 c74 (.A(net6),
    .B(net861),
    .X(net12));
 sky130_fd_sc_hd__sdfbbn_1 c740 (.CLK_N(clknet_4_7_0_clk),
    .D(net1049),
    .RESET_B(net526),
    .SCD(net594),
    .SCE(net596),
    .SET_B(net681),
    .Q(net608));
 sky130_fd_sc_hd__or4bb_1 c741 (.A(net608),
    .B(net943),
    .C_N(net602),
    .D_N(net460),
    .X(net609));
 sky130_fd_sc_hd__sdfbbn_1 c742 (.CLK_N(clknet_4_7_0_clk),
    .D(net526),
    .RESET_B(net460),
    .SCD(net943),
    .SCE(net601),
    .SET_B(net681),
    .Q(net610));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net610),
    .A1(net460),
    .A2(net601),
    .A3(net599),
    .S0(net995),
    .S1(net809),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net545),
    .A1(net579),
    .A2(net602),
    .A3(net594),
    .S0(net951),
    .S1(net717),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net612),
    .A1(net603),
    .A2(net602),
    .A3(net943),
    .S0(net954),
    .S1(net545),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net943),
    .A1(net962),
    .A2(net971),
    .A3(net800),
    .S0(net805),
    .S1(net808),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net481),
    .A1(net594),
    .A2(net478),
    .A3(net943),
    .S0(net807),
    .S1(net812),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net577),
    .A1(clknet_1_1__leaf_net595),
    .A2(net575),
    .A3(net985),
    .S0(net874),
    .S1(net719),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net527),
    .A1(net530),
    .A2(net848),
    .A3(clknet_1_0__leaf_net595),
    .S0(net798),
    .S1(clknet_1_0__leaf_net806),
    .X(net617));
 sky130_fd_sc_hd__and2_4 c75 (.A(net10),
    .B(net12),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net500),
    .A1(net481),
    .A2(clknet_1_0__leaf_net595),
    .A3(net713),
    .S0(net783),
    .S1(clknet_1_1__leaf_net806),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(clknet_1_1__leaf_net482),
    .A1(net481),
    .A2(clknet_1_0__leaf_net595),
    .A3(net527),
    .S0(net783),
    .S1(net796),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net223),
    .A1(net527),
    .A2(net575),
    .A3(net963),
    .S0(net805),
    .S1(net813),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net874),
    .A1(net574),
    .A2(net832),
    .A3(net868),
    .S0(net798),
    .S1(net813),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net874),
    .A1(clknet_1_1__leaf_net707),
    .A2(net721),
    .A3(net796),
    .S0(net798),
    .S1(clknet_1_1__leaf_net806),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net530),
    .A1(clknet_1_0__leaf_net622),
    .A2(net575),
    .A3(net720),
    .S0(net971),
    .S1(clknet_1_1__leaf_net806),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net585),
    .A1(net499),
    .A2(net530),
    .A3(net733),
    .S1(net796),
    .X(net742));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net954),
    .A1(net989),
    .A2(net741),
    .A3(net796),
    .S0(net798),
    .S1(net813),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net621),
    .A1(net575),
    .A2(clknet_1_1__leaf_net595),
    .A3(net805),
    .S0(clknet_1_1__leaf_net806),
    .S1(net813),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(clknet_1_1__leaf_net595),
    .A1(net986),
    .A2(net623),
    .A3(clknet_1_1__leaf_net622),
    .S0(net782),
    .S1(net813),
    .X(net627));
 sky130_fd_sc_hd__and3_1 c76 (.A(net858),
    .B(net10),
    .C(net830),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net13),
    .A1(clknet_1_1__leaf_net595),
    .A2(net527),
    .A3(net625),
    .S0(net971),
    .S1(net813),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(clknet_1_1__leaf_net595),
    .A1(net735),
    .A2(net796),
    .A3(net805),
    .S0(net811),
    .S1(net814),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net625),
    .A1(net703),
    .A2(net905),
    .A3(net810),
    .S0(net813),
    .S1(net814),
    .X(net630));
 sky130_fd_sc_hd__and3_1 c77 (.A(net12),
    .B(net9),
    .C(net10),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c78 (.A(net849),
    .B(net854),
    .X(net16));
 sky130_fd_sc_hd__a2111o_1 c79 (.A1(net858),
    .A2(net10),
    .B1(net13),
    .C1(net879),
    .D1(net16),
    .X(net17));
 sky130_fd_sc_hd__and2_0 c80 (.A(net11),
    .B(net15),
    .X(net18));
 sky130_fd_sc_hd__and2_1 c81 (.A(net830),
    .B(net13),
    .X(net19));
 sky130_fd_sc_hd__mux4_2 c82 (.A0(net12),
    .A1(net18),
    .A2(net11),
    .A3(net2),
    .S0(net865),
    .S1(net15),
    .X(net20));
 sky130_fd_sc_hd__and2_1 c83 (.A(net18),
    .B(net20),
    .X(net21));
 sky130_fd_sc_hd__and2_1 c84 (.A(net21),
    .B(net17),
    .X(net22));
 sky130_fd_sc_hd__or4bb_4 c85 (.A(net15),
    .B(net16),
    .C_N(net21),
    .D_N(net825),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net16),
    .A1(net11),
    .A2(net21),
    .A3(net23),
    .S0(net873),
    .S1(net22),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net4),
    .A1(net864),
    .A2(net7),
    .A3(net24),
    .S0(net847),
    .S1(net23),
    .X(net918));
 sky130_fd_sc_hd__and2_1 c88 (.A(net8),
    .B(net841),
    .X(net25));
 sky130_fd_sc_hd__and2_1 c89 (.A(net9),
    .B(net22),
    .X(net26));
 sky130_fd_sc_hd__and2_1 c90 (.A(net841),
    .B(net874),
    .X(net27));
 sky130_fd_sc_hd__and2_1 c91 (.A(net21),
    .B(net26),
    .X(net28));
 sky130_fd_sc_hd__and3_2 c92 (.A(net4),
    .B(net28),
    .C(net9),
    .X(net29));
 sky130_fd_sc_hd__and3_1 c93 (.A(net959),
    .B(net28),
    .C(net25),
    .X(net30));
 sky130_fd_sc_hd__and2_2 c94 (.A(net832),
    .B(net30),
    .X(net31));
 sky130_fd_sc_hd__and2_1 c95 (.A(net25),
    .B(net28),
    .X(net32));
 sky130_fd_sc_hd__or4bb_4 c96 (.A(net870),
    .B(net14),
    .C_N(net4),
    .D_N(net950),
    .X(net33));
 sky130_fd_sc_hd__and2_0 c97 (.A(net14),
    .B(net27),
    .X(net34));
 sky130_fd_sc_hd__and2_0 c98 (.A(net28),
    .B(net1),
    .X(net35));
 sky130_fd_sc_hd__and2_2 c99 (.A(net6),
    .B(net32),
    .X(net36));
 sky130_fd_sc_hd__mux4_1 merge763 (.A0(net963),
    .A1(net411),
    .A2(clknet_1_0__leaf_net477),
    .A3(net883),
    .S0(net223),
    .S1(net555),
    .X(net631));
 sky130_fd_sc_hd__a2111o_1 merge764 (.A1(net103),
    .A2(net848),
    .B1(net966),
    .C1(net211),
    .D1(net114),
    .X(net632));
 sky130_fd_sc_hd__a2111o_1 merge765 (.A1(net108),
    .A2(net873),
    .B1(net107),
    .C1(net105),
    .D1(net95),
    .X(net633));
 sky130_fd_sc_hd__or4bb_1 merge766 (.A(net41),
    .B(net54),
    .C_N(net745),
    .D_N(net747),
    .X(net634));
 sky130_fd_sc_hd__sedfxtp_1 merge767 (.CLK(clknet_4_9_0_clk),
    .D(net363),
    .DE(net956),
    .SCD(net343),
    .SCE(net737),
    .Q(net635));
 sky130_fd_sc_hd__mux4_1 merge768 (.A0(net538),
    .A1(net867),
    .A2(net947),
    .A3(net546),
    .S0(net85),
    .S1(net787),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 merge769 (.A(net700),
    .X(net637));
 sky130_fd_sc_hd__sdfbbp_1 merge770 (.CLK(clknet_4_0_0_clk),
    .D(net84),
    .RESET_B(net952),
    .SCD(net945),
    .SCE(net212),
    .SET_B(net1040),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__or4bb_1 merge771 (.A(net23),
    .B(net124),
    .C_N(net92),
    .D_N(net871),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 merge772 (.A(net819),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net37),
    .A1(net45),
    .A2(net152),
    .A3(net60),
    .S0(net976),
    .S1(net41),
    .X(net642));
 sky130_fd_sc_hd__or4bb_1 merge774 (.A(net103),
    .B(net216),
    .C_N(net212),
    .D_N(net728),
    .X(net643));
 sky130_fd_sc_hd__or4bb_1 merge775 (.A(net295),
    .B(net313),
    .C_N(net202),
    .D_N(net835),
    .X(net644));
 sky130_fd_sc_hd__sedfxtp_1 merge776 (.CLK(clknet_4_8_0_clk),
    .D(net145),
    .DE(net981),
    .SCD(net92),
    .SCE(net33),
    .Q(net645));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net97),
    .A1(net296),
    .A2(net946),
    .A3(net338),
    .S0(net944),
    .S1(net874),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net869),
    .A1(net262),
    .A2(net967),
    .A3(clknet_1_1__leaf_net154),
    .S0(net269),
    .S1(net940),
    .X(net647));
 sky130_fd_sc_hd__a2111o_1 merge779 (.A1(net524),
    .A2(net539),
    .B1(net527),
    .C1(net533),
    .D1(net680),
    .X(net648));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net105),
    .A1(net133),
    .A2(net137),
    .A3(net834),
    .S0(net98),
    .S1(net202),
    .X(net649));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net313),
    .A1(clknet_1_0__leaf_net482),
    .A2(clknet_1_1__leaf_net480),
    .A3(net587),
    .S0(clknet_1_1__leaf_net708),
    .S1(net801),
    .X(net650));
 sky130_fd_sc_hd__or4bb_1 merge782 (.A(net198),
    .B(net295),
    .C_N(net303),
    .D_N(net294),
    .X(net651));
 sky130_fd_sc_hd__sdfrbp_1 merge783 (.CLK(clknet_4_8_0_clk),
    .D(net145),
    .RESET_B(net5),
    .SCD(net45),
    .SCE(clknet_1_0__leaf_net754),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__a2111o_1 merge784 (.A1(net916),
    .A2(net294),
    .B1(net195),
    .C1(net198),
    .D1(net973),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net543),
    .A1(net538),
    .A2(net573),
    .A3(net944),
    .S0(net205),
    .S1(net225),
    .X(net655));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net438),
    .A1(net313),
    .A2(net311),
    .A3(net337),
    .S0(clknet_1_0__leaf_net771),
    .S1(net787),
    .X(net656));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net327),
    .A1(net556),
    .A2(net573),
    .A3(net530),
    .S0(clknet_1_1__leaf_net771),
    .S1(net772),
    .X(net657));
 sky130_fd_sc_hd__a2111o_1 merge788 (.A1(net184),
    .A2(net198),
    .B1(net203),
    .C1(net217),
    .D1(net212),
    .X(net658));
 sky130_fd_sc_hd__sdfbbn_1 merge789 (.CLK_N(clknet_4_10_0_clk),
    .D(net166),
    .RESET_B(clknet_1_1__leaf_net930),
    .SCD(net172),
    .SCE(net911),
    .SET_B(net1029),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net58),
    .A1(net45),
    .A2(net55),
    .A3(net170),
    .S0(net911),
    .S1(net926),
    .X(net661));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net96),
    .A1(net269),
    .A2(net227),
    .A3(net982),
    .S0(net271),
    .S1(net270),
    .X(net662));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net108),
    .A1(net954),
    .A2(net109),
    .A3(net224),
    .S0(net236),
    .S1(net211),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net235),
    .A1(net236),
    .A2(net963),
    .A3(net242),
    .S0(net877),
    .S1(net237),
    .X(net664));
 sky130_fd_sc_hd__a2111o_1 merge794 (.A1(net440),
    .A2(net960),
    .B1(net947),
    .C1(net417),
    .D1(net962),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net155),
    .A1(net42),
    .A2(net32),
    .A3(net41),
    .S0(net903),
    .S1(net967),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net7),
    .A1(net133),
    .A2(net937),
    .A3(net915),
    .S0(net949),
    .S1(net958),
    .X(net667));
 sky130_fd_sc_hd__a2111o_1 merge797 (.A1(net171),
    .A2(net170),
    .B1(net45),
    .C1(net903),
    .D1(net750),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net311),
    .A1(net961),
    .A2(net454),
    .A3(net523),
    .S0(net679),
    .S1(net804),
    .X(net669));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net171),
    .A1(net64),
    .A2(net923),
    .A3(net847),
    .S0(net1051),
    .S1(net937),
    .X(net670));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net295),
    .A1(net973),
    .A2(net198),
    .A3(net828),
    .S0(net229),
    .S1(net202),
    .X(net671));
 sky130_fd_sc_hd__dfrbp_1 merge801 (.CLK(clknet_4_12_0_clk),
    .D(net383),
    .RESET_B(net390),
    .Q(net672),
    .Q_N(net914));
 sky130_fd_sc_hd__dfrbp_1 merge802 (.CLK(clknet_4_6_0_clk),
    .D(net494),
    .RESET_B(net491),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net201),
    .B(net658),
    .X(net675));
 sky130_fd_sc_hd__and2_4 merge804 (.A(net570),
    .B(net571),
    .X(net676));
 sky130_fd_sc_hd__and2_0 merge805 (.A(net630),
    .B(net616),
    .X(net677));
 sky130_fd_sc_hd__and2_0 merge806 (.A(net275),
    .B(net288),
    .X(net678));
 sky130_fd_sc_hd__dfrtn_1 merge807 (.CLK_N(clknet_4_4_0_clk),
    .D(net426),
    .Q(net427));
 sky130_fd_sc_hd__dfrtp_1 merge808 (.CLK(clknet_4_10_0_clk),
    .D(net51),
    .RESET_B(net63),
    .Q(net888));
 sky130_fd_sc_hd__dfrtp_1 merge809 (.CLK(clknet_4_5_0_clk),
    .D(net541),
    .RESET_B(net544),
    .Q(net680));
 sky130_fd_sc_hd__dfrtp_1 merge810 (.CLK(clknet_4_7_0_clk),
    .D(net597),
    .RESET_B(net598),
    .Q(net681));
 sky130_fd_sc_hd__dfsbp_1 merge811 (.CLK(clknet_4_6_0_clk),
    .D(net453),
    .SET_B(net455),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__dfsbp_1 merge812 (.CLK(clknet_4_9_0_clk),
    .D(net266),
    .SET_B(net247),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__dfstp_1 merge813 (.CLK(clknet_4_2_0_clk),
    .D(net632),
    .SET_B(net664),
    .Q(net686));
 sky130_fd_sc_hd__and2_0 merge814 (.A(net358),
    .B(net360),
    .X(net687));
 sky130_fd_sc_hd__dfstp_1 merge815 (.CLK(clknet_4_0_0_clk),
    .D(net104),
    .Q(net106));
 sky130_fd_sc_hd__dfstp_1 merge816 (.CLK(clknet_4_1_0_clk),
    .D(net431),
    .SET_B(net439),
    .Q(net689));
 sky130_fd_sc_hd__dlrbn_1 merge817 (.D(net380),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net382),
    .Q(net907),
    .Q_N(net690));
 sky130_fd_sc_hd__and2_0 merge818 (.A(net178),
    .B(net180),
    .X(net691));
 sky130_fd_sc_hd__and2_0 merge819 (.A(net643),
    .B(net213),
    .X(net692));
 sky130_fd_sc_hd__dlrbn_1 merge820 (.GATE_N(clknet_4_11_0_clk),
    .RESET_B(net292),
    .Q(net891),
    .Q_N(net293));
 sky130_fd_sc_hd__dlrbp_1 merge821 (.D(net503),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net505),
    .Q(net941),
    .Q_N(net694));
 sky130_fd_sc_hd__and2_0 merge822 (.A(net127),
    .B(net633),
    .X(net695));
 sky130_fd_sc_hd__dlrbp_1 merge823 (.D(net164),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net157),
    .Q(net900),
    .Q_N(net696));
 sky130_fd_sc_hd__dlrtn_1 merge824 (.D(net318),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net319),
    .Q(net697));
 sky130_fd_sc_hd__and2_0 merge825 (.A(net139),
    .B(net147),
    .X(net698));
 sky130_fd_sc_hd__dlrtn_1 merge826 (.D(net566),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net550),
    .Q(net699));
 sky130_fd_sc_hd__dlrtn_1 merge827 (.D(net651),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net654),
    .Q(net700));
 sky130_fd_sc_hd__dlrtp_1 merge828 (.D(net43),
    .GATE(clknet_4_8_0_clk),
    .Q(net44));
 sky130_fd_sc_hd__dlrtp_1 merge829 (.D(net644),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net648),
    .Q(net702));
 sky130_fd_sc_hd__dlrtp_1 merge830 (.D(net512),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net629),
    .Q(net703));
 sky130_fd_sc_hd__edfxbp_1 merge831 (.CLK(clknet_4_1_0_clk),
    .DE(net687),
    .Q(net361),
    .Q_N(net704));
 sky130_fd_sc_hd__edfxtp_1 merge832 (.CLK(clknet_4_12_0_clk),
    .D(net341),
    .DE(net381),
    .Q(net706));
 sky130_fd_sc_hd__sdlclkp_1 merge833 (.CLK(clknet_4_6_0_clk),
    .GATE(net677),
    .SCE(net461),
    .GCLK(net707));
 sky130_fd_sc_hd__sdlclkp_2 merge834 (.CLK(clknet_4_6_0_clk),
    .GATE(net470),
    .SCE(net591),
    .GCLK(net708));
 sky130_fd_sc_hd__and2_0 merge835 (.A(net391),
    .B(net521),
    .X(net709));
 sky130_fd_sc_hd__sdlclkp_4 merge836 (.CLK(clknet_4_15_0_clk),
    .GATE(net471),
    .SCE(net518),
    .GCLK(net710));
 sky130_fd_sc_hd__dfrbp_1 merge837 (.CLK(clknet_4_0_0_clk),
    .D(net671),
    .RESET_B(net320),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dfrbp_1 merge838 (.CLK(clknet_4_7_0_clk),
    .D(net604),
    .RESET_B(net615),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__and2_0 merge839 (.A(net181),
    .B(net397),
    .X(net715));
 sky130_fd_sc_hd__dfrtn_1 merge840 (.CLK_N(clknet_4_3_0_clk),
    .D(net472),
    .RESET_B(net334),
    .Q(net716));
 sky130_fd_sc_hd__dfrtp_1 merge841 (.CLK(clknet_4_13_0_clk),
    .D(net517),
    .RESET_B(net627),
    .Q(net905));
 sky130_fd_sc_hd__dfrtp_1 merge842 (.CLK(clknet_4_7_0_clk),
    .D(net609),
    .RESET_B(net590),
    .Q(net717));
 sky130_fd_sc_hd__and2_0 merge843 (.A(net640),
    .B(net261),
    .X(net718));
 sky130_fd_sc_hd__dfrtp_1 merge844 (.CLK(clknet_4_12_0_clk),
    .D(net509),
    .RESET_B(net398),
    .Q(net719));
 sky130_fd_sc_hd__dfsbp_1 merge845 (.CLK(clknet_4_13_0_clk),
    .D(net617),
    .SET_B(net618),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dfsbp_1 merge846 (.CLK(clknet_4_2_0_clk),
    .D(net663),
    .SET_B(net695),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dfstp_1 merge847 (.CLK(clknet_4_11_0_clk),
    .D(net678),
    .SET_B(net662),
    .Q(net724));
 sky130_fd_sc_hd__and2_0 merge848 (.A(net200),
    .B(net675),
    .X(net725));
 sky130_fd_sc_hd__dfstp_1 merge849 (.CLK(clknet_4_9_0_clk),
    .D(net647),
    .SET_B(net715),
    .Q(net726));
 sky130_fd_sc_hd__dfstp_1 merge850 (.CLK(clknet_4_10_0_clk),
    .D(net634),
    .SET_B(net670),
    .Q(net727));
 sky130_fd_sc_hd__dlrbn_2 merge851 (.D(net725),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net692),
    .Q(net729),
    .Q_N(net728));
 sky130_fd_sc_hd__dlrbn_1 merge852 (.D(net691),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net649),
    .Q(net898),
    .Q_N(net730));
 sky130_fd_sc_hd__dlrbp_1 merge853 (.D(net405),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net401),
    .Q(net917),
    .Q_N(net731));
 sky130_fd_sc_hd__dlrbp_1 merge854 (.D(net676),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net450),
    .Q(net733),
    .Q_N(net732));
 sky130_fd_sc_hd__dlrtn_2 merge855 (.D(net253),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net709),
    .Q(net734));
 sky130_fd_sc_hd__dlrtn_1 merge856 (.D(net600),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net626),
    .Q(net735));
 sky130_fd_sc_hd__and2_0 merge857 (.A(net667),
    .B(net698),
    .X(net736));
 sky130_fd_sc_hd__dlrtn_2 merge858 (.D(net718),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net736),
    .Q(net737));
 sky130_fd_sc_hd__dlrtp_1 merge859 (.D(net646),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net321),
    .Q(net738));
 sky130_fd_sc_hd__dlrtp_1 merge860 (.D(net669),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net665),
    .Q(net739));
 sky130_fd_sc_hd__dlrtp_1 merge861 (.D(net326),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net636),
    .Q(net740));
 sky130_fd_sc_hd__edfxbp_1 merge862 (.CLK(clknet_4_15_0_clk),
    .D(net620),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__edfxtp_1 merge863 (.CLK(clknet_4_10_0_clk),
    .D(net159),
    .DE(net668),
    .Q(net743));
 sky130_fd_sc_hd__sdlclkp_1 merge864 (.CLK(clknet_4_5_0_clk),
    .GATE(net565),
    .SCE(net655),
    .GCLK(net744));
 sky130_fd_sc_hd__dfxbp_1 s865 (.CLK(clknet_4_10_0_clk),
    .D(net40),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__dfxbp_1 s866 (.CLK(clknet_4_10_0_clk),
    .D(net46),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dfxtp_2 s867 (.CLK(clknet_4_10_0_clk),
    .D(net57),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_1 s868 (.CLK(clknet_4_10_0_clk),
    .D(net59),
    .Q(net750));
 sky130_fd_sc_hd__dfxtp_2 s869 (.CLK(clknet_4_8_0_clk),
    .D(net146),
    .Q(net751));
 sky130_fd_sc_hd__dlclkp_1 s870 (.CLK(clknet_4_8_0_clk),
    .GATE(net150),
    .GCLK(net752));
 sky130_fd_sc_hd__dlclkp_2 s871 (.CLK(clknet_4_8_0_clk),
    .GATE(net153),
    .GCLK(net753));
 sky130_fd_sc_hd__dlclkp_4 s872 (.CLK(clknet_4_8_0_clk),
    .GATE(net160),
    .GCLK(net754));
 sky130_fd_sc_hd__dlxbn_1 s873 (.D(net167),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net935),
    .Q_N(net755));
 sky130_fd_sc_hd__dlxbn_1 s874 (.D(net176),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net757),
    .Q_N(net756));
 sky130_fd_sc_hd__dlxbp_1 s875 (.D(net244),
    .GATE(clknet_4_2_0_clk),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__dlxtn_2 s876 (.D(net265),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net940));
 sky130_fd_sc_hd__dlxtn_1 s877 (.D(net274),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net760));
 sky130_fd_sc_hd__dlxtn_1 s878 (.D(net277),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net761));
 sky130_fd_sc_hd__dlxtp_1 s879 (.D(net281),
    .GATE(clknet_4_11_0_clk),
    .Q(net762));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s880 (.D(net283),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net929));
 sky130_fd_sc_hd__dfxbp_1 s881 (.CLK(clknet_4_11_0_clk),
    .D(net287),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dfxbp_1 s882 (.CLK(clknet_4_11_0_clk),
    .D(net289),
    .Q(net766),
    .Q_N(net765));
 sky130_fd_sc_hd__dfxtp_4 s883 (.CLK(clknet_4_11_0_clk),
    .D(net290),
    .Q(net767));
 sky130_fd_sc_hd__dfxtp_1 s884 (.CLK(clknet_4_11_0_clk),
    .D(net291),
    .Q(net931));
 sky130_fd_sc_hd__dfxtp_2 s885 (.CLK(clknet_4_1_0_clk),
    .D(net310),
    .Q(net768));
 sky130_fd_sc_hd__dlclkp_1 s886 (.CLK(clknet_4_0_0_clk),
    .GATE(net329),
    .GCLK(net769));
 sky130_fd_sc_hd__dlclkp_2 s887 (.CLK(clknet_4_2_0_clk),
    .GATE(net330),
    .GCLK(net770));
 sky130_fd_sc_hd__dlclkp_4 s888 (.CLK(clknet_4_1_0_clk),
    .GATE(net331),
    .GCLK(net771));
 sky130_fd_sc_hd__dlxbn_1 s889 (.D(net335),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__dlxbn_1 s890 (.D(net354),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net775),
    .Q_N(net774));
 sky130_fd_sc_hd__dlxbp_1 s891 (.D(net355),
    .GATE(clknet_4_3_0_clk),
    .Q(net777),
    .Q_N(net776));
 sky130_fd_sc_hd__dlxtn_2 s892 (.D(net370),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net901));
 sky130_fd_sc_hd__dlxtn_1 s893 (.D(net371),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net778));
 sky130_fd_sc_hd__dlxtn_1 s894 (.D(net379),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net779));
 sky130_fd_sc_hd__dlxtp_1 s895 (.D(net384),
    .GATE(clknet_4_14_0_clk),
    .Q(net780));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s896 (.D(net387),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net781));
 sky130_fd_sc_hd__dfxbp_1 s897 (.CLK(clknet_4_13_0_clk),
    .D(net407),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dfxbp_1 s898 (.CLK(clknet_4_4_0_clk),
    .D(net424),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dfxtp_1 s899 (.CLK(clknet_4_4_0_clk),
    .D(net428),
    .Q(net786));
 sky130_fd_sc_hd__dfxtp_2 s900 (.CLK(clknet_4_1_0_clk),
    .D(net447),
    .Q(net787));
 sky130_fd_sc_hd__dfxtp_1 s901 (.CLK(clknet_4_4_0_clk),
    .D(net449),
    .Q(net788));
 sky130_fd_sc_hd__dlclkp_1 s902 (.CLK(clknet_4_6_0_clk),
    .GATE(net462),
    .GCLK(net884));
 sky130_fd_sc_hd__dlclkp_2 s903 (.CLK(clknet_4_6_0_clk),
    .GATE(net465),
    .GCLK(net789));
 sky130_fd_sc_hd__dlclkp_4 s904 (.CLK(clknet_4_12_0_clk),
    .GATE(net492),
    .GCLK(net892));
 sky130_fd_sc_hd__dlxbn_1 s905 (.D(net506),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net896),
    .Q_N(net790));
 sky130_fd_sc_hd__dlxbn_1 s906 (.D(net508),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net897),
    .Q_N(net791));
 sky130_fd_sc_hd__dlxbp_1 s907 (.D(net511),
    .GATE(clknet_4_12_0_clk),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__dlxtn_2 s908 (.D(net513),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net794));
 sky130_fd_sc_hd__dlxtn_1 s909 (.D(net514),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net795));
 sky130_fd_sc_hd__dlxtn_1 s910 (.D(net516),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net796));
 sky130_fd_sc_hd__dlxtp_1 s911 (.D(net519),
    .GATE(clknet_4_15_0_clk),
    .Q(net797));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s912 (.D(net522),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net798));
 sky130_fd_sc_hd__dfxbp_1 s913 (.CLK(clknet_4_7_0_clk),
    .D(net551),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dfxbp_1 s914 (.CLK(clknet_4_5_0_clk),
    .D(net563),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dfxtp_1 s915 (.CLK(clknet_4_5_0_clk),
    .D(net564),
    .Q(net803));
 sky130_fd_sc_hd__dfxtp_1 s916 (.CLK(clknet_4_5_0_clk),
    .D(net568),
    .Q(net804));
 sky130_fd_sc_hd__dfxtp_2 s917 (.CLK(clknet_4_7_0_clk),
    .D(net588),
    .Q(net805));
 sky130_fd_sc_hd__dlclkp_1 s918 (.CLK(clknet_4_7_0_clk),
    .GATE(net589),
    .GCLK(net806));
 sky130_fd_sc_hd__dlclkp_2 s919 (.CLK(clknet_4_7_0_clk),
    .GATE(net605),
    .GCLK(net807));
 sky130_fd_sc_hd__dlclkp_4 s920 (.CLK(clknet_4_13_0_clk),
    .GATE(net606),
    .GCLK(net808));
 sky130_fd_sc_hd__dlxbn_1 s921 (.D(net607),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dlxbn_1 s922 (.D(net611),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net810));
 sky130_fd_sc_hd__dlxbp_1 s923 (.D(net613),
    .GATE(clknet_4_13_0_clk),
    .Q(net811));
 sky130_fd_sc_hd__dlxtn_1 s924 (.D(net614),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net812));
 sky130_fd_sc_hd__dlxtn_2 s925 (.D(net619),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net813));
 sky130_fd_sc_hd__dlxtn_1 s926 (.D(net628),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net814));
 sky130_fd_sc_hd__dlxtp_1 s927 (.D(net631),
    .GATE(clknet_4_4_0_clk),
    .Q(net815));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s928 (.D(net642),
    .SLEEP_B(clknet_4_10_0_clk),
    .Q(net816));
 sky130_fd_sc_hd__dfxbp_1 s929 (.CLK(clknet_4_6_0_clk),
    .D(net650),
    .Q(net818),
    .Q_N(net817));
 sky130_fd_sc_hd__dfxbp_1 s930 (.CLK(clknet_4_4_0_clk),
    .D(net656),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__dfxtp_1 s931 (.CLK(clknet_4_6_0_clk),
    .D(net657),
    .Q(net821));
 sky130_fd_sc_hd__dfxtp_1 s932 (.CLK(clknet_4_10_0_clk),
    .D(net661),
    .Q(net822));
 sky130_fd_sc_hd__dfxtp_1 s933 (.CLK(clknet_4_10_0_clk),
    .D(net666),
    .Q(net823));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in0),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net825));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net827));
 sky130_fd_sc_hd__buf_6 input7 (.A(in14),
    .X(net828));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(in15),
    .X(net829));
 sky130_fd_sc_hd__buf_1 input9 (.A(in16),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net831));
 sky130_fd_sc_hd__buf_12 input11 (.A(in18),
    .X(net832));
 sky130_fd_sc_hd__buf_1 input12 (.A(in19),
    .X(net833));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net834));
 sky130_fd_sc_hd__buf_8 input14 (.A(in20),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in21),
    .X(net836));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(in22),
    .X(net837));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input21 (.A(in27),
    .X(net842));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input25 (.A(in30),
    .X(net846));
 sky130_fd_sc_hd__buf_2 input26 (.A(in31),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(in32),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input29 (.A(in34),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input31 (.A(in36),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input32 (.A(in37),
    .X(net853));
 sky130_fd_sc_hd__buf_1 input33 (.A(in38),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net855));
 sky130_fd_sc_hd__buf_1 input35 (.A(in4),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in40),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in41),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in42),
    .X(net859));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net860));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(in44),
    .X(net861));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(in45),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net863));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(in48),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(in5),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(in50),
    .X(net868));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net869));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net870));
 sky130_fd_sc_hd__buf_2 input50 (.A(in53),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in54),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(in55),
    .X(net873));
 sky130_fd_sc_hd__buf_4 input53 (.A(in56),
    .X(net874));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net875));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net876));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net877));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net878));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in61),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(in7),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in8),
    .X(net882));
 sky130_fd_sc_hd__buf_4 input62 (.A(in9),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(clknet_1_1__leaf_net884),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net885),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output65 (.A(net886),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(clknet_1_1__leaf_net887),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output67 (.A(net888),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(clknet_1_1__leaf_net889),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net890),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output70 (.A(net891),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(clknet_1_1__leaf_net892),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output72 (.A(net960),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output73 (.A(net894),
    .X(out19));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net895),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output75 (.A(net896),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output76 (.A(net897),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output77 (.A(net898),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output78 (.A(net899),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output79 (.A(net900),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output80 (.A(net901),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output81 (.A(net902),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output82 (.A(net903),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output83 (.A(net904),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net905),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output85 (.A(net906),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output86 (.A(net907),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output87 (.A(net908),
    .X(out32));
 sky130_fd_sc_hd__buf_2 output88 (.A(net909),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net910),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output90 (.A(net911),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output91 (.A(net912),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output92 (.A(net913),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output93 (.A(net914),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output94 (.A(net915),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output95 (.A(net916),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output96 (.A(net917),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net978),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(clknet_1_1__leaf_net919),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net920),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output100 (.A(net921),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net922),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output102 (.A(net923),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output103 (.A(net924),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output104 (.A(net925),
    .X(out48));
 sky130_fd_sc_hd__buf_2 output105 (.A(net926),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output106 (.A(net927),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output107 (.A(net928),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output108 (.A(net929),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(clknet_1_0__leaf_net930),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output110 (.A(net931),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output111 (.A(net932),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output112 (.A(net933),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output113 (.A(net934),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output114 (.A(net935),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output115 (.A(net936),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output116 (.A(net937),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output117 (.A(net952),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output118 (.A(net939),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output119 (.A(net940),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output120 (.A(net941),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net942),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net599),
    .X(net943));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net327),
    .X(net944));
 sky130_fd_sc_hd__buf_2 fanout124 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net948),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net948),
    .X(net947));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net314),
    .X(net948));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(net249),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net31),
    .X(net950));
 sky130_fd_sc_hd__buf_12 fanout130 (.A(net561),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net938),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net123),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net101),
    .X(net954));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net460),
    .X(net955));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net364),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net225),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net29),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net893),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net429),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net885),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net233),
    .X(net963));
 sky130_fd_sc_hd__buf_12 fanout143 (.A(net894),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net968),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net116),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net435),
    .X(net969));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net255),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net788),
    .X(net971));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net187),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(net187),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net806 (.A(net806),
    .X(clknet_0_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_0__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net806 (.A(clknet_0_net806),
    .X(clknet_1_1__leaf_net806));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net622 (.A(net622),
    .X(clknet_0_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_0__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net622 (.A(clknet_0_net622),
    .X(clknet_1_1__leaf_net622));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net708 (.A(net708),
    .X(clknet_0_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_0__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_1__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net892 (.A(net892),
    .X(clknet_0_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_0__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net892 (.A(clknet_0_net892),
    .X(clknet_1_1__leaf_net892));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net789 (.A(net789),
    .X(clknet_0_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_0__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net789 (.A(clknet_0_net789),
    .X(clknet_1_1__leaf_net789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net480 (.A(net480),
    .X(clknet_0_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net480 (.A(clknet_0_net480),
    .X(clknet_1_0__leaf_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net480 (.A(clknet_0_net480),
    .X(clknet_1_1__leaf_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net482 (.A(net482),
    .X(clknet_0_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_0__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net482 (.A(clknet_0_net482),
    .X(clknet_1_1__leaf_net482));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net477 (.A(net477),
    .X(clknet_0_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_0__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_1__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net771 (.A(net771),
    .X(clknet_0_net771));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net771 (.A(clknet_0_net771),
    .X(clknet_1_0__leaf_net771));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net771 (.A(clknet_0_net771),
    .X(clknet_1_1__leaf_net771));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net770 (.A(net770),
    .X(clknet_0_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net770 (.A(clknet_0_net770),
    .X(clknet_1_1__leaf_net770));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net507 (.A(net507),
    .X(clknet_0_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_0__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net507 (.A(clknet_0_net507),
    .X(clknet_1_1__leaf_net507));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net769 (.A(net769),
    .X(clknet_0_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_0__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net769 (.A(clknet_0_net769),
    .X(clknet_1_1__leaf_net769));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net754 (.A(net754),
    .X(clknet_0_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net754 (.A(clknet_0_net754),
    .X(clknet_1_0__leaf_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net754 (.A(clknet_0_net754),
    .X(clknet_1_1__leaf_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net168 (.A(net168),
    .X(clknet_0_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_0__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net168 (.A(clknet_0_net168),
    .X(clknet_1_1__leaf_net168));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net753 (.A(net753),
    .X(clknet_0_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_0__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_1__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net930 (.A(net930),
    .X(clknet_0_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_0__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net930 (.A(clknet_0_net930),
    .X(clknet_1_1__leaf_net930));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net154 (.A(net154),
    .X(clknet_0_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_0__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net154 (.A(clknet_0_net154),
    .X(clknet_1_1__leaf_net154));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net752 (.A(net752),
    .X(clknet_0_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_0__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_1__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net887 (.A(net887),
    .X(clknet_0_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net887 (.A(clknet_0_net887),
    .X(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net919 (.A(net919),
    .X(clknet_0_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_1__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net889 (.A(net889),
    .X(clknet_0_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net744 (.A(net744),
    .X(clknet_0_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_0__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net744 (.A(clknet_0_net744),
    .X(clknet_1_1__leaf_net744));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net344 (.A(net344),
    .X(clknet_0_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_0__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net344 (.A(clknet_0_net344),
    .X(clknet_1_1__leaf_net344));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net359 (.A(net359),
    .X(clknet_0_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_0__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net359 (.A(clknet_0_net359),
    .X(clknet_1_1__leaf_net359));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net373 (.A(net373),
    .X(clknet_0_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_0__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net373 (.A(clknet_0_net373),
    .X(clknet_1_1__leaf_net373));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net376 (.A(net376),
    .X(clknet_0_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_0__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net376 (.A(clknet_0_net376),
    .X(clknet_1_1__leaf_net376));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net710 (.A(net710),
    .X(clknet_0_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_0__leaf_net710));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net710 (.A(clknet_0_net710),
    .X(clknet_1_1__leaf_net710));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net824),
    .A1(net826),
    .A2(net70),
    .A3(net68),
    .S0(net964),
    .S1(net624),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net918),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net918),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net976),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net976),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net24),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net979),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net979),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net979),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net979),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net0),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net984),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net985),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net67),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net67),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer16 (.A(net988),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net894),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net337),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net81),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net97),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net308),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net1002),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net97),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net964),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 clone25 (.A(net894),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net20),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net999),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net1000),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1018),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net702),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net1064),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net489),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net448),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net672),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net767),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net787),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net487),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net781),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net731),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net55),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net267),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net711),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net697),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net474),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net328),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net680),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net908),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net356),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net931),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net716),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net579),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net859),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net60),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net817),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net766),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net796),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net762),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net802),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net396),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net764),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net804),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net760),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net759),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net746),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net388),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net749),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net429),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net748),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net888),
    .X(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_D (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SCE (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_D1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_Q (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_SCE (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_C_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_D_N (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_D1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_D_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_C (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_D_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_C_N (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_D_N (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCE (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_D1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_RESET_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_C_N (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_D_N (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_S0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCE (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_D1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SET_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_D (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_C (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q_N (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_C_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_C1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SCD (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_D1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_C1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCD (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A0 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCE (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_C1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_D (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCE (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_SCD (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_Q (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_Q (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_RESET_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_C (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_C_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_D_N (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SET_B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_SCE (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_C1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_S0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SET_B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C_N (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_C (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_C1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_B1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_C_N (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCE (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_SCD (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_RESET_B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_C (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_Q_N (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_RESET_B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_D_N (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_GATE (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_D (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_RESET_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_X (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCD (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_C_N (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_C (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A0 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_RESET_B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCD (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_Q (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_D1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_B (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_X (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer15_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_D1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_RESET_B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_D (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold75_A (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_Q_N (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_D_N (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_D1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_Q (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_D_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_D1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_Q (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_SCE (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_SCE (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D_N (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_C (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold60_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_Q (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SET_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_C1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_C1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_C (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net770_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GCLK (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_Q_N (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold81_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_Q (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_C (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_Q_N (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_D1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_Q (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_D (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_D1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCD (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_C_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_C1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_C1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_D1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_S1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_D_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_C (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_C (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_C (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_C (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_C1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_D_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_C (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SCE (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold77_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A0 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_D_N (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_C (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_C_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_SET_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_C_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_D_N (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_B1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A2 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_D_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_SCD (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_C (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_C (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_C1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_C1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net887_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone25_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_SET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_X (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_RESET_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_RESET_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_SCE (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_D_N (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_SCE (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_Q (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCD (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_Q (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_SCE (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_C1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_SCD (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_Q (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_SCD (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_SCE (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCD (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_RESET_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A2 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_Q (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_C (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_C (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_SET_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_Q (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_SCE (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_D (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_D_N (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_SCD (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_RESET_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_C1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_D_N (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_D1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_SCD (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_SET_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_RESET_B (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SET_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SET_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_RESET_B (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_C_N (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCD (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_SCE (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_D1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_C1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SCD (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_SCD (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCD (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_D_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_D1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_C_N (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_SET_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_RESET_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_SCE (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_D1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_D1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_C (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_C1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_D_N (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_C1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_C_N (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_D1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_C_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_D1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_D_N (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_RESET_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_C1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_C1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_D_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_D_N (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_SCE (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_C1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_C_N (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_D1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_C (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_SCE (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_D (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_B1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_C_N (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_D_N (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_C (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_D1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_D1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_C (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_D1 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_C_N (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S0 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_D_N (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_C (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_D1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_C1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_D_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_C (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_SLEEP_B (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_D1 (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SET_B (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_D1 (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_D1 (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D_N (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net884_X (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_C1 (.DIODE(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net884_X (.DIODE(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net770_X (.DIODE(clknet_1_0__leaf_net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S1 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net887_X (.DIODE(clknet_1_0__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_C1 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_C1 (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net887_X (.DIODE(clknet_1_1__leaf_net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B (.DIODE(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net372_X (.DIODE(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone1_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_S0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_C1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_C_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SCE (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCE (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone25_X (.DIODE(net998));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net824),
    .A1(net826),
    .A2(net70),
    .A3(net68),
    .S0(net964),
    .S1(net624),
    .X(net1003));
 sky130_fd_sc_hd__a2111o_1 clone3 (.A1(net17),
    .A2(net113),
    .B1(net131),
    .C1(net125),
    .D1(net92),
    .X(net1004));
 sky130_fd_sc_hd__and3_1 clone4 (.A(net69),
    .B(net66),
    .C(net70),
    .X(net1005));
 sky130_fd_sc_hd__and3_1 clone5 (.A(net67),
    .B(net881),
    .C(net832),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net77),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net1007),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net1007),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1007),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net77),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net1011),
    .X(net1012));
 sky130_fd_sc_hd__mux4_1 clone35 (.A0(net1020),
    .A1(net336),
    .A2(net301),
    .A3(net332),
    .S0(net738),
    .S1(net773),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net1),
    .X(net1014));
 sky130_fd_sc_hd__and3_1 clone37 (.A(net66),
    .B(net65),
    .C(net826),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(in18),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net561),
    .X(net1018));
 sky130_fd_sc_hd__or4bb_1 clone41 (.A(net91),
    .B(net90),
    .C_N(net852),
    .D_N(net859),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net308),
    .X(net1020));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
