module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net668;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net905;
 wire clknet_1_0__leaf_net905;
 wire clknet_1_1__leaf_net905;
 wire clknet_0_net738;
 wire clknet_1_0__leaf_net738;
 wire clknet_1_1__leaf_net738;
 wire clknet_0_net276;
 wire clknet_1_0__leaf_net276;
 wire clknet_1_1__leaf_net276;
 wire clknet_0_net279;
 wire clknet_1_0__leaf_net279;
 wire clknet_1_1__leaf_net279;
 wire clknet_0_net408;
 wire clknet_1_0__leaf_net408;
 wire clknet_1_1__leaf_net408;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net502;
 wire clknet_1_0__leaf_net502;
 wire clknet_1_1__leaf_net502;
 wire clknet_0_net964;
 wire clknet_1_0__leaf_net964;
 wire clknet_1_1__leaf_net964;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net412;
 wire clknet_1_0__leaf_net412;
 wire clknet_1_1__leaf_net412;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net410;
 wire clknet_1_0__leaf_net410;
 wire clknet_1_1__leaf_net410;
 wire clknet_0_net270;
 wire clknet_1_0__leaf_net270;
 wire clknet_1_1__leaf_net270;
 wire clknet_0_net273;
 wire clknet_1_0__leaf_net273;
 wire clknet_1_1__leaf_net273;
 wire clknet_0_net730;
 wire clknet_1_0__leaf_net730;
 wire clknet_1_1__leaf_net730;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net814;
 wire clknet_1_0__leaf_net814;
 wire clknet_1_1__leaf_net814;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net304;
 wire clknet_1_0__leaf_net304;
 wire clknet_1_1__leaf_net304;
 wire clknet_0_net473;
 wire clknet_1_0__leaf_net473;
 wire clknet_1_1__leaf_net473;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net459;
 wire clknet_1_0__leaf_net459;
 wire clknet_1_1__leaf_net459;
 wire clknet_0_net464;
 wire clknet_1_0__leaf_net464;
 wire clknet_1_1__leaf_net464;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net587;
 wire clknet_1_0__leaf_net587;
 wire clknet_1_1__leaf_net587;
 wire clknet_0_net582;
 wire clknet_1_0__leaf_net582;
 wire clknet_1_1__leaf_net582;
 wire clknet_0_net695;
 wire clknet_1_0__leaf_net695;
 wire clknet_1_1__leaf_net695;
 wire clknet_0_net816;
 wire clknet_1_0__leaf_net816;
 wire clknet_1_1__leaf_net816;
 wire clknet_0_net333;
 wire clknet_1_0__leaf_net333;
 wire clknet_1_1__leaf_net333;
 wire clknet_0_net300;
 wire clknet_1_0__leaf_net300;
 wire clknet_1_1__leaf_net300;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire clknet_0_net963;
 wire clknet_1_0__leaf_net963;
 wire clknet_1_1__leaf_net963;
 wire clknet_0_net869;
 wire clknet_1_0__leaf_net869;
 wire clknet_1_1__leaf_net869;
 wire clknet_0_net498;
 wire clknet_1_0__leaf_net498;
 wire clknet_1_1__leaf_net498;
 wire clknet_0_net314;
 wire clknet_1_0__leaf_net314;
 wire clknet_1_1__leaf_net314;
 wire clknet_0_net287;
 wire clknet_1_0__leaf_net287;
 wire clknet_1_1__leaf_net287;
 wire clknet_0_net313;
 wire clknet_1_0__leaf_net313;
 wire clknet_1_1__leaf_net313;
 wire clknet_0_net309;
 wire clknet_1_0__leaf_net309;
 wire clknet_1_1__leaf_net309;
 wire clknet_0_net290;
 wire clknet_1_0__leaf_net290;
 wire clknet_1_1__leaf_net290;
 wire clknet_0_net903;
 wire clknet_1_0__leaf_net903;
 wire clknet_1_1__leaf_net903;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net586;
 wire clknet_1_0__leaf_net586;
 wire clknet_1_1__leaf_net586;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net886;
 wire clknet_1_0__leaf_net886;
 wire clknet_1_1__leaf_net886;
 wire clknet_0_net885;
 wire clknet_1_0__leaf_net885;
 wire clknet_1_1__leaf_net885;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net680;
 wire clknet_1_0__leaf_net680;
 wire clknet_1_1__leaf_net680;
 wire clknet_0_net679;
 wire clknet_1_0__leaf_net679;
 wire clknet_1_1__leaf_net679;
 wire clknet_0_net681;
 wire clknet_1_0__leaf_net681;
 wire clknet_1_1__leaf_net681;
 wire clknet_0_net851;
 wire clknet_1_0__leaf_net851;
 wire clknet_1_1__leaf_net851;
 wire clknet_0_net850;
 wire clknet_1_0__leaf_net850;
 wire clknet_1_1__leaf_net850;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net830;
 wire clknet_1_0__leaf_net830;
 wire clknet_1_1__leaf_net830;
 wire clknet_0_net219;
 wire clknet_1_0__leaf_net219;
 wire clknet_1_1__leaf_net219;
 wire clknet_0_net230;
 wire clknet_1_0__leaf_net230;
 wire clknet_1_1__leaf_net230;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net218;
 wire clknet_1_0__leaf_net218;
 wire clknet_1_1__leaf_net218;
 wire clknet_0_net217;
 wire clknet_1_0__leaf_net217;
 wire clknet_1_1__leaf_net217;
 wire clknet_0_net216;
 wire clknet_1_0__leaf_net216;
 wire clknet_1_1__leaf_net216;
 wire clknet_0_net828;
 wire clknet_1_0__leaf_net828;
 wire clknet_1_1__leaf_net828;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;

 sky130_fd_sc_hd__clkbuf_2 c100 (.A(net810),
    .X(net73));
 sky130_fd_sc_hd__xnor2_1 c101 (.A(net65),
    .B(net73),
    .Y(net74));
 sky130_fd_sc_hd__buf_1 c102 (.A(net756),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net74),
    .A1(net47),
    .A2(net66),
    .A3(net73),
    .S0(net68),
    .S1(net795),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 c104 (.A(net911),
    .X(net77));
 sky130_fd_sc_hd__a21bo_2 c105 (.A1(net73),
    .A2(net3),
    .B1_N(net972),
    .X(net78));
 sky130_fd_sc_hd__sdfrbp_1 c106 (.CLK(clknet_4_13_0_clk),
    .D(net72),
    .RESET_B(net69),
    .SCD(net73),
    .SCE(net972),
    .Q(net80),
    .Q_N(net79));
 sky130_fd_sc_hd__mux4_1 c107 (.A0(net71),
    .A1(net74),
    .A2(net973),
    .A3(net79),
    .S0(net73),
    .S1(net795),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net69),
    .A1(net77),
    .A2(net73),
    .A3(net982),
    .S0(net1038),
    .S1(net972),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net77),
    .A1(net78),
    .A2(net82),
    .A3(net73),
    .S0(net41),
    .S1(net65),
    .X(net83));
 sky130_fd_sc_hd__xnor2_1 c110 (.A(net982),
    .B(net19),
    .Y(net84));
 sky130_fd_sc_hd__xnor2_2 c111 (.A(net44),
    .B(net48),
    .Y(net85));
 sky130_fd_sc_hd__a41o_1 c112 (.A1(net72),
    .A2(net64),
    .A3(net975),
    .A4(net810),
    .B1(net1063),
    .X(net86));
 sky130_fd_sc_hd__xnor2_4 c113 (.A(net51),
    .B(net1027),
    .Y(net87));
 sky130_fd_sc_hd__a31o_1 c114 (.A1(net33),
    .A2(net59),
    .A3(net981),
    .B1(net973),
    .X(net88));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net88),
    .B(net973),
    .Y(net89));
 sky130_fd_sc_hd__dfbbn_1 c116 (.CLK_N(clknet_4_13_0_clk),
    .D(net89),
    .RESET_B(net44),
    .SET_B(net827),
    .Q(net91),
    .Q_N(net90));
 sky130_fd_sc_hd__a21bo_1 c117 (.A1(net64),
    .A2(net967),
    .B1_N(net87),
    .X(net92));
 sky130_fd_sc_hd__buf_2 c118 (.A(net1072),
    .X(net93));
 sky130_fd_sc_hd__buf_1 c119 (.A(net908),
    .X(net94));
 sky130_fd_sc_hd__xnor2_2 c120 (.A(net94),
    .B(net87),
    .Y(net95));
 sky130_fd_sc_hd__xnor2_2 c121 (.A(net91),
    .B(net93),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_1 c122 (.A(net59),
    .B(net94),
    .Y(net97));
 sky130_fd_sc_hd__sdfrbp_2 c123 (.CLK(clknet_4_15_0_clk),
    .D(net95),
    .RESET_B(net85),
    .SCD(net90),
    .SCE(net975),
    .Q(net99),
    .Q_N(net98));
 sky130_fd_sc_hd__clkbuf_1 c124 (.A(net1072),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 c125 (.A(net910),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 c126 (.A0(net87),
    .A1(net90),
    .A2(net95),
    .A3(net98),
    .S0(net93),
    .S1(net1070),
    .X(net102));
 sky130_fd_sc_hd__a21bo_1 c127 (.A1(net100),
    .A2(net87),
    .B1_N(net975),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net48),
    .A1(net989),
    .A2(net92),
    .A3(net91),
    .S0(net103),
    .S1(net981),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net103),
    .A1(net99),
    .A2(net974),
    .A3(net45),
    .S0(net1063),
    .S1(clknet_1_1__leaf_net828),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c130 (.A0(net103),
    .A1(net95),
    .A2(net99),
    .A3(net64),
    .S0(net788),
    .S1(clknet_1_1__leaf_net828),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net85),
    .A1(net974),
    .A2(net103),
    .A3(net810),
    .S0(net950),
    .S1(net829),
    .X(net107));
 sky130_fd_sc_hd__buf_4 c132 (.A(net939),
    .X(net108));
 sky130_fd_sc_hd__buf_2 c133 (.A(net928),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 c134 (.A(net923),
    .X(net110));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net925),
    .B(net921),
    .Y(net111));
 sky130_fd_sc_hd__clkbuf_4 c136 (.A(net931),
    .X(net112));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net929),
    .B(net1008),
    .Y(net113));
 sky130_fd_sc_hd__xnor2_4 c138 (.A(net941),
    .B(net1008),
    .Y(net114));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net924),
    .B(net923),
    .Y(net115));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net114),
    .B(net115),
    .Y(net116));
 sky130_fd_sc_hd__xnor2_4 c141 (.A(net939),
    .B(net116),
    .Y(net117));
 sky130_fd_sc_hd__xnor2_2 c142 (.A(net113),
    .B(net934),
    .Y(net118));
 sky130_fd_sc_hd__xnor2_4 c143 (.A(net1003),
    .B(net112),
    .Y(net119));
 sky130_fd_sc_hd__xnor2_4 c144 (.A(net108),
    .B(net113),
    .Y(net120));
 sky130_fd_sc_hd__a21bo_4 c145 (.A1(net118),
    .A2(net1003),
    .B1_N(net127),
    .X(net121));
 sky130_fd_sc_hd__xnor2_4 c146 (.A(net121),
    .B(net1014),
    .Y(net122));
 sky130_fd_sc_hd__a21bo_4 c147 (.A1(net112),
    .A2(net120),
    .B1_N(net121),
    .X(net123));
 sky130_fd_sc_hd__xnor2_4 c148 (.A(net121),
    .B(net123),
    .Y(net965));
 sky130_fd_sc_hd__a21bo_2 c149 (.A1(net116),
    .A2(net119),
    .B1_N(net123),
    .X(net124));
 sky130_fd_sc_hd__xnor2_4 c150 (.A(net1003),
    .B(net121),
    .Y(net125));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net109),
    .A1(net124),
    .A2(net123),
    .A3(net125),
    .S0(net117),
    .S1(net120),
    .X(net126));
 sky130_fd_sc_hd__xnor2_4 c152 (.A(net122),
    .B(net991),
    .Y(net959));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net120),
    .A1(net113),
    .A2(net117),
    .A3(net118),
    .S0(net115),
    .S1(net1008),
    .X(net127));
 sky130_fd_sc_hd__xnor2_4 c154 (.A(net124),
    .B(net125),
    .Y(net128));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net986),
    .B(net8),
    .Y(net129));
 sky130_fd_sc_hd__xnor2_2 c156 (.A(net12),
    .B(net668),
    .Y(net130));
 sky130_fd_sc_hd__xnor2_4 c157 (.A(net129),
    .B(net989),
    .Y(net968));
 sky130_fd_sc_hd__xnor2_2 c158 (.A(net5),
    .B(net18),
    .Y(net131));
 sky130_fd_sc_hd__xnor2_4 c159 (.A(net112),
    .B(net128),
    .Y(net957));
 sky130_fd_sc_hd__xnor2_2 c160 (.A(net15),
    .B(net129),
    .Y(net132));
 sky130_fd_sc_hd__xnor2_4 c161 (.A(net12),
    .B(net995),
    .Y(net133));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net928),
    .B(net923),
    .Y(net134));
 sky130_fd_sc_hd__mux4_2 c163 (.A0(net921),
    .A1(net15),
    .A2(net968),
    .A3(net131),
    .S0(net13),
    .S1(net985),
    .X(net135));
 sky130_fd_sc_hd__xnor2_2 c164 (.A(net923),
    .B(net15),
    .Y(net136));
 sky130_fd_sc_hd__xnor2_2 c165 (.A(net132),
    .B(net968),
    .Y(net137));
 sky130_fd_sc_hd__xnor2_2 c166 (.A(net129),
    .B(net136),
    .Y(net138));
 sky130_fd_sc_hd__xnor2_1 c167 (.A(net933),
    .B(net985),
    .Y(net139));
 sky130_fd_sc_hd__xnor2_1 c168 (.A(net941),
    .B(net977),
    .Y(net951));
 sky130_fd_sc_hd__xnor2_2 c169 (.A(net131),
    .B(net977),
    .Y(net140));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net136),
    .A1(net124),
    .A2(net128),
    .A3(net135),
    .S0(net133),
    .S1(net977),
    .X(net141));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net141),
    .A1(net135),
    .A2(net132),
    .A3(net977),
    .S0(net133),
    .S1(net139),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net142),
    .A1(net985),
    .A2(net141),
    .A3(net938),
    .S0(net136),
    .S1(net977),
    .X(net143));
 sky130_fd_sc_hd__buf_1 c173 (.A(net821),
    .X(net144));
 sky130_fd_sc_hd__xnor2_4 c174 (.A(net140),
    .B(net1022),
    .Y(net145));
 sky130_fd_sc_hd__clkbuf_1 c175 (.A(net821),
    .X(net146));
 sky130_fd_sc_hd__a21bo_1 c176 (.A1(net122),
    .A2(net145),
    .B1_N(net8),
    .X(net147));
 sky130_fd_sc_hd__a21bo_1 c177 (.A1(net21),
    .A2(net22),
    .B1_N(net1006),
    .X(net148));
 sky130_fd_sc_hd__xnor2_2 c178 (.A(net118),
    .B(net18),
    .Y(net149));
 sky130_fd_sc_hd__xnor2_2 c179 (.A(net34),
    .B(net145),
    .Y(net150));
 sky130_fd_sc_hd__xnor2_4 c180 (.A(net122),
    .B(net35),
    .Y(net151));
 sky130_fd_sc_hd__xnor2_4 c181 (.A(net995),
    .B(net151),
    .Y(net152));
 sky130_fd_sc_hd__buf_1 c182 (.A(net790),
    .X(net153));
 sky130_fd_sc_hd__xnor2_1 c183 (.A(net152),
    .B(net149),
    .Y(net154));
 sky130_fd_sc_hd__xnor2_1 c184 (.A(net38),
    .B(net927),
    .Y(net155));
 sky130_fd_sc_hd__a31o_1 c185 (.A1(net139),
    .A2(net150),
    .A3(net30),
    .B1(net152),
    .X(net156));
 sky130_fd_sc_hd__xnor2_1 c186 (.A(net21),
    .B(net821),
    .Y(net157));
 sky130_fd_sc_hd__clkbuf_4 c187 (.A(net755),
    .X(net158));
 sky130_fd_sc_hd__xnor2_2 c188 (.A(net151),
    .B(net821),
    .Y(net159));
 sky130_fd_sc_hd__xnor2_2 c189 (.A(net153),
    .B(net8),
    .Y(net160));
 sky130_fd_sc_hd__clkbuf_1 c190 (.A(net790),
    .X(net161));
 sky130_fd_sc_hd__buf_2 c191 (.A(net764),
    .X(net162));
 sky130_fd_sc_hd__xnor2_2 c192 (.A(net1085),
    .B(net162),
    .Y(net163));
 sky130_fd_sc_hd__a21bo_1 c193 (.A1(net161),
    .A2(net163),
    .B1_N(net26),
    .X(net164));
 sky130_fd_sc_hd__sdfrtn_1 c194 (.CLK_N(clknet_4_7_0_clk),
    .D(net164),
    .RESET_B(net163),
    .SCD(net1002),
    .SCE(net30),
    .Q(net165));
 sky130_fd_sc_hd__a21bo_1 c195 (.A1(net161),
    .A2(net1002),
    .B1_N(net165),
    .X(net166));
 sky130_fd_sc_hd__a41o_1 c196 (.A1(net148),
    .A2(net164),
    .A3(net133),
    .A4(net166),
    .B1(net668),
    .X(net167));
 sky130_fd_sc_hd__a41o_4 c197 (.A1(net166),
    .A2(net162),
    .A3(net8),
    .A4(net1002),
    .B1(net791),
    .X(net168));
 sky130_fd_sc_hd__xnor2_1 c198 (.A(net55),
    .B(net165),
    .Y(net169));
 sky130_fd_sc_hd__a21bo_2 c199 (.A1(net31),
    .A2(net148),
    .B1_N(net989),
    .X(net170));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net1086),
    .A2(net170),
    .B1_N(net55),
    .X(net171));
 sky130_fd_sc_hd__a41o_1 c201 (.A1(net154),
    .A2(net55),
    .A3(net948),
    .A4(net1002),
    .B1(net51),
    .X(net172));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net49),
    .A2(net1011),
    .B1_N(net821),
    .X(net173));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net921),
    .A2(net160),
    .B1_N(net111),
    .X(net174));
 sky130_fd_sc_hd__a21bo_1 c204 (.A1(net171),
    .A2(net165),
    .B1_N(net1086),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c205 (.A1(net153),
    .A2(net169),
    .B1_N(net813),
    .X(net176));
 sky130_fd_sc_hd__buf_2 c206 (.A(net813),
    .X(net177));
 sky130_fd_sc_hd__xnor2_4 c207 (.A(net158),
    .B(net813),
    .Y(net178));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(net49),
    .A2(net111),
    .B1_N(net986),
    .X(net179));
 sky130_fd_sc_hd__a21bo_2 c209 (.A1(net986),
    .A2(net174),
    .B1_N(net176),
    .X(net180));
 sky130_fd_sc_hd__xnor2_1 c210 (.A(net32),
    .B(net813),
    .Y(net181));
 sky130_fd_sc_hd__a31o_1 c211 (.A1(net50),
    .A2(net181),
    .A3(net923),
    .B1(net31),
    .X(net182));
 sky130_fd_sc_hd__a31o_1 c212 (.A1(net181),
    .A2(net1086),
    .A3(net177),
    .B1(net170),
    .X(net183));
 sky130_fd_sc_hd__a21bo_1 c213 (.A1(net174),
    .A2(net178),
    .B1_N(net182),
    .X(net184));
 sky130_fd_sc_hd__a21bo_1 c214 (.A1(net184),
    .A2(net170),
    .B1_N(net813),
    .X(net185));
 sky130_fd_sc_hd__buf_2 c215 (.A(net813),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net182),
    .A1(net157),
    .A2(net986),
    .A3(net186),
    .S0(net50),
    .S1(net821),
    .X(net187));
 sky130_fd_sc_hd__a21bo_1 c217 (.A1(net187),
    .A2(net149),
    .B1_N(net170),
    .X(net188));
 sky130_fd_sc_hd__a21bo_1 c218 (.A1(net185),
    .A2(net186),
    .B1_N(net188),
    .X(net189));
 sky130_fd_sc_hd__a41o_1 c219 (.A1(net176),
    .A2(net1006),
    .A3(net188),
    .A4(net182),
    .B1(net180),
    .X(net190));
 sky130_fd_sc_hd__a21bo_2 c220 (.A1(net149),
    .A2(net45),
    .B1_N(net972),
    .X(net191));
 sky130_fd_sc_hd__a21bo_1 c221 (.A1(net995),
    .A2(net186),
    .B1_N(net78),
    .X(net192));
 sky130_fd_sc_hd__a21bo_1 c222 (.A1(net51),
    .A2(net170),
    .B1_N(net1006),
    .X(net193));
 sky130_fd_sc_hd__a21bo_1 c223 (.A1(net165),
    .A2(net173),
    .B1_N(net180),
    .X(net194));
 sky130_fd_sc_hd__buf_1 c224 (.A(net786),
    .X(net195));
 sky130_fd_sc_hd__xnor2_1 c225 (.A(net32),
    .B(net178),
    .Y(net196));
 sky130_fd_sc_hd__a31o_1 c226 (.A1(net196),
    .A2(net173),
    .A3(net191),
    .B1(net825),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 c227 (.A(net786),
    .X(net198));
 sky130_fd_sc_hd__a21bo_1 c228 (.A1(net26),
    .A2(net196),
    .B1_N(net198),
    .X(net199));
 sky130_fd_sc_hd__a31o_1 c229 (.A1(net173),
    .A2(net54),
    .A3(net191),
    .B1(net198),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net148),
    .A1(net191),
    .A2(net1012),
    .A3(net198),
    .S0(net193),
    .S1(net795),
    .X(net201));
 sky130_fd_sc_hd__sdfbbn_1 c231 (.CLK_N(clknet_4_12_0_clk),
    .D(net192),
    .RESET_B(net46),
    .SCD(net972),
    .SCE(net173),
    .SET_B(net795),
    .Q(net203),
    .Q_N(net202));
 sky130_fd_sc_hd__clkbuf_1 c232 (.A(net907),
    .X(net204));
 sky130_fd_sc_hd__a41o_1 c233 (.A1(net193),
    .A2(net202),
    .A3(net178),
    .A4(net957),
    .B1(net972),
    .X(net205));
 sky130_fd_sc_hd__xnor2_1 c234 (.A(net170),
    .B(net826),
    .Y(net206));
 sky130_fd_sc_hd__buf_6 c235 (.A(net906),
    .X(net207));
 sky130_fd_sc_hd__sdfbbn_2 c236 (.CLK_N(clknet_4_13_0_clk),
    .D(net1006),
    .RESET_B(net1052),
    .SCD(net51),
    .SCE(net1043),
    .SET_B(net192),
    .Q(net209),
    .Q_N(net208));
 sky130_fd_sc_hd__a21bo_4 c237 (.A1(net135),
    .A2(net204),
    .B1_N(net207),
    .X(net210));
 sky130_fd_sc_hd__mux4_1 c238 (.A0(net200),
    .A1(net203),
    .A2(net205),
    .A3(net1043),
    .S0(net13),
    .S1(net972),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net205),
    .A1(net198),
    .A2(net206),
    .A3(net23),
    .S0(net1042),
    .S1(net974),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c240 (.A0(net204),
    .A1(net957),
    .A2(net207),
    .A3(net192),
    .S0(net786),
    .S1(net831),
    .X(net213));
 sky130_fd_sc_hd__sdfbbp_1 c241 (.CLK(clknet_4_12_0_clk),
    .D(net201),
    .RESET_B(net160),
    .SCD(net208),
    .SCE(net832),
    .SET_B(net834),
    .Q(net215),
    .Q_N(net214));
 sky130_fd_sc_hd__a21bo_4 c242 (.A1(net210),
    .A2(net162),
    .B1_N(net93),
    .X(net947));
 sky130_fd_sc_hd__a21bo_1 c243 (.A1(net96),
    .A2(net206),
    .B1_N(clknet_1_0__leaf_net830),
    .X(net216));
 sky130_fd_sc_hd__a31o_1 c244 (.A1(net947),
    .A2(net162),
    .A3(net974),
    .B1(clknet_1_1__leaf_net830),
    .X(net217));
 sky130_fd_sc_hd__a31o_1 c245 (.A1(net80),
    .A2(net1030),
    .A3(net826),
    .B1(clknet_1_1__leaf_net830),
    .X(net218));
 sky130_fd_sc_hd__a21bo_1 c246 (.A1(net974),
    .A2(net826),
    .B1_N(clknet_1_0__leaf_net830),
    .X(net219));
 sky130_fd_sc_hd__a31o_1 c247 (.A1(clknet_1_1__leaf_net216),
    .A2(net198),
    .A3(clknet_1_0__leaf_net219),
    .B1(net974),
    .X(net220));
 sky130_fd_sc_hd__sdfrtp_1 c248 (.CLK(clknet_4_13_0_clk),
    .D(net975),
    .RESET_B(net85),
    .SCD(net194),
    .SCE(clknet_1_0__leaf_net830),
    .Q(net221));
 sky130_fd_sc_hd__sdfbbn_1 c249 (.CLK_N(clknet_4_15_0_clk),
    .D(net85),
    .RESET_B(clknet_1_1__leaf_net220),
    .SCD(net1005),
    .SCE(clknet_1_1__leaf_net828),
    .SET_B(clknet_1_1__leaf_net830),
    .Q(net223),
    .Q_N(net222));
 sky130_fd_sc_hd__xnor2_4 c25 (.A(net939),
    .B(net937),
    .Y(net0));
 sky130_fd_sc_hd__sdfbbn_1 c250 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_0__leaf_net220),
    .RESET_B(net210),
    .SCD(net96),
    .SCE(net974),
    .SET_B(net791),
    .Q(net966),
    .Q_N(net224));
 sky130_fd_sc_hd__sdfrtp_2 c251 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net219),
    .RESET_B(clknet_1_0__leaf_net220),
    .SCD(net1005),
    .SCE(net96),
    .Q(net225));
 sky130_fd_sc_hd__a41o_1 c252 (.A1(net194),
    .A2(net198),
    .A3(net225),
    .A4(net974),
    .B1(net101),
    .X(net958));
 sky130_fd_sc_hd__a31o_1 c253 (.A1(net225),
    .A2(net194),
    .A3(net1005),
    .B1(net795),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(net206),
    .A1(net958),
    .A2(net79),
    .A3(net208),
    .S0(net1005),
    .S1(net98),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net45),
    .A1(net227),
    .A2(net80),
    .A3(net226),
    .S0(net974),
    .S1(net168),
    .X(net228));
 sky130_fd_sc_hd__a41o_1 c256 (.A1(net198),
    .A2(net1065),
    .A3(net226),
    .A4(net1005),
    .B1(net194),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(net225),
    .A1(net226),
    .A2(net96),
    .A3(clknet_1_0__leaf_net219),
    .S0(net974),
    .S1(clknet_1_0__leaf_net216),
    .X(net230));
 sky130_fd_sc_hd__sdfbbp_1 c258 (.CLK(clknet_4_15_0_clk),
    .D(net226),
    .RESET_B(net1005),
    .SCD(clknet_1_0__leaf_net230),
    .SCE(net1065),
    .SET_B(net227),
    .Q(net232),
    .Q_N(net231));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net101),
    .A1(net958),
    .A2(clknet_1_1__leaf_net219),
    .A3(clknet_1_1__leaf_net220),
    .S0(clknet_1_0__leaf_net230),
    .S1(net222),
    .X(net233));
 sky130_fd_sc_hd__xnor2_4 c26 (.A(net935),
    .B(net933),
    .Y(net1));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(clknet_1_1__leaf_net230),
    .A1(net232),
    .A2(net85),
    .A3(net225),
    .S0(net1005),
    .S1(clknet_1_1__leaf_net830),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(clknet_1_1__leaf_net217),
    .A1(clknet_1_0__leaf_net230),
    .A2(net222),
    .A3(net98),
    .S0(net823),
    .S1(net825),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net221),
    .A1(clknet_1_1__leaf_net230),
    .A2(net231),
    .A3(net803),
    .S0(net822),
    .S1(net837),
    .X(net236));
 sky130_fd_sc_hd__sdfbbn_1 c263 (.CLK_N(clknet_4_15_0_clk),
    .D(net1041),
    .RESET_B(clknet_1_1__leaf_net230),
    .SCD(net804),
    .SCE(net1073),
    .SET_B(net1053),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net668),
    .B(net1007),
    .Y(net239));
 sky130_fd_sc_hd__clkbuf_2 c265 (.A(net924),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 c266 (.A(net933),
    .X(net241));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net1009),
    .B(net108),
    .Y(net242));
 sky130_fd_sc_hd__xnor2_2 c268 (.A(net240),
    .B(net1007),
    .Y(net243));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net242),
    .B(net1001),
    .Y(net244));
 sky130_fd_sc_hd__xnor2_4 c27 (.A(net929),
    .B(net0),
    .Y(net2));
 sky130_fd_sc_hd__a31o_4 c270 (.A1(net1007),
    .A2(net240),
    .A3(net126),
    .B1(net110),
    .X(net245));
 sky130_fd_sc_hd__xnor2_1 c271 (.A(net240),
    .B(net924),
    .Y(net246));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net239),
    .B(net242),
    .Y(net247));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net119),
    .B(net241),
    .Y(net248));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net244),
    .B(net126),
    .Y(net249));
 sky130_fd_sc_hd__xnor2_4 c275 (.A(net926),
    .B(net245),
    .Y(net250));
 sky130_fd_sc_hd__xnor2_2 c276 (.A(net242),
    .B(net978),
    .Y(net251));
 sky130_fd_sc_hd__xnor2_2 c277 (.A(net119),
    .B(net110),
    .Y(net252));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net247),
    .B(net927),
    .Y(net253));
 sky130_fd_sc_hd__xnor2_1 c279 (.A(net253),
    .B(net247),
    .Y(net254));
 sky130_fd_sc_hd__xnor2_4 c28 (.A(net943),
    .B(net937),
    .Y(net3));
 sky130_fd_sc_hd__xnor2_4 c280 (.A(net253),
    .B(net932),
    .Y(net255));
 sky130_fd_sc_hd__xnor2_4 c281 (.A(net252),
    .B(net984),
    .Y(net256));
 sky130_fd_sc_hd__xnor2_2 c282 (.A(net244),
    .B(net255),
    .Y(net257));
 sky130_fd_sc_hd__xnor2_4 c283 (.A(net978),
    .B(net245),
    .Y(net258));
 sky130_fd_sc_hd__xnor2_4 c284 (.A(net251),
    .B(net256),
    .Y(net259));
 sky130_fd_sc_hd__xnor2_4 c285 (.A(net259),
    .B(net258),
    .Y(net260));
 sky130_fd_sc_hd__xnor2_2 c286 (.A(net120),
    .B(net977),
    .Y(net261));
 sky130_fd_sc_hd__xnor2_1 c287 (.A(net1),
    .B(net243),
    .Y(net262));
 sky130_fd_sc_hd__xnor2_2 c288 (.A(net991),
    .B(net243),
    .Y(net263));
 sky130_fd_sc_hd__xnor2_1 c289 (.A(net254),
    .B(net1010),
    .Y(net264));
 sky130_fd_sc_hd__a21bo_4 c29 (.A1(net938),
    .A2(net930),
    .B1_N(net1),
    .X(net4));
 sky130_fd_sc_hd__a21bo_1 c290 (.A1(net146),
    .A2(net256),
    .B1_N(net989),
    .X(net265));
 sky130_fd_sc_hd__xnor2_4 c291 (.A(net991),
    .B(net263),
    .Y(net266));
 sky130_fd_sc_hd__xnor2_4 c292 (.A(net239),
    .B(net668),
    .Y(net267));
 sky130_fd_sc_hd__xnor2_2 c293 (.A(net265),
    .B(net145),
    .Y(net268));
 sky130_fd_sc_hd__xnor2_4 c294 (.A(net4),
    .B(net267),
    .Y(net269));
 sky130_fd_sc_hd__buf_1 c295 (.A(clknet_1_1__leaf_net738),
    .X(net270));
 sky130_fd_sc_hd__xnor2_2 c296 (.A(net265),
    .B(net668),
    .Y(net271));
 sky130_fd_sc_hd__xnor2_1 c297 (.A(net13),
    .B(net1),
    .Y(net272));
 sky130_fd_sc_hd__xnor2_1 c298 (.A(net271),
    .B(clknet_1_1__leaf_net270),
    .Y(net273));
 sky130_fd_sc_hd__clkbuf_2 c299 (.A(net762),
    .X(net274));
 sky130_fd_sc_hd__xnor2_4 c30 (.A(net1),
    .B(net943),
    .Y(net5));
 sky130_fd_sc_hd__a41o_1 c300 (.A1(clknet_1_0__leaf_net270),
    .A2(net264),
    .A3(net254),
    .A4(net142),
    .B1(net994),
    .X(net275));
 sky130_fd_sc_hd__buf_1 c301 (.A(clknet_1_0__leaf_net738),
    .X(net276));
 sky130_fd_sc_hd__xnor2_4 c302 (.A(net15),
    .B(net274),
    .Y(net277));
 sky130_fd_sc_hd__a31o_1 c303 (.A1(net272),
    .A2(net994),
    .A3(net984),
    .B1(net145),
    .X(net278));
 sky130_fd_sc_hd__a41o_1 c304 (.A1(clknet_1_0__leaf_net276),
    .A2(net138),
    .A3(net134),
    .A4(net668),
    .B1(net266),
    .X(net279));
 sky130_fd_sc_hd__a31o_1 c305 (.A1(net275),
    .A2(net272),
    .A3(clknet_1_1__leaf_net276),
    .B1(net971),
    .X(net280));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net263),
    .A2(net278),
    .A3(net138),
    .A4(net277),
    .X(net281));
 sky130_fd_sc_hd__a41o_2 c307 (.A1(net8),
    .A2(net146),
    .A3(net269),
    .A4(net258),
    .B1(net787),
    .X(net282));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net264),
    .B(net978),
    .Y(net283));
 sky130_fd_sc_hd__xnor2_4 c309 (.A(net33),
    .B(net787),
    .Y(net284));
 sky130_fd_sc_hd__xnor2_4 c31 (.A(net5),
    .B(net0),
    .Y(net6));
 sky130_fd_sc_hd__xnor2_2 c310 (.A(net36),
    .B(net137),
    .Y(net285));
 sky130_fd_sc_hd__buf_1 c311 (.A(net913),
    .X(net286));
 sky130_fd_sc_hd__buf_1 c312 (.A(clknet_1_1__leaf_net730),
    .X(net287));
 sky130_fd_sc_hd__xnor2_2 c313 (.A(net277),
    .B(net787),
    .Y(net288));
 sky130_fd_sc_hd__buf_1 c314 (.A(clknet_1_0__leaf_net730),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net277),
    .A1(net145),
    .A2(clknet_1_0__leaf_net287),
    .A3(net152),
    .S0(net668),
    .S1(net133),
    .X(net290));
 sky130_fd_sc_hd__xnor2_1 c316 (.A(net289),
    .B(net37),
    .Y(net291));
 sky130_fd_sc_hd__clkbuf_2 c317 (.A(net763),
    .X(net292));
 sky130_fd_sc_hd__a21bo_1 c318 (.A1(net145),
    .A2(net286),
    .B1_N(net668),
    .X(net293));
 sky130_fd_sc_hd__xnor2_1 c319 (.A(net283),
    .B(net168),
    .Y(net294));
 sky130_fd_sc_hd__a21bo_1 c32 (.A1(net4),
    .A2(net5),
    .B1_N(net928),
    .X(net7));
 sky130_fd_sc_hd__xnor2_1 c320 (.A(clknet_1_0__leaf_net291),
    .B(net288),
    .Y(net295));
 sky130_fd_sc_hd__buf_1 c321 (.A(clknet_1_1__leaf_net814),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net147),
    .A1(clknet_1_1__leaf_net291),
    .A2(net292),
    .A3(net288),
    .S0(clknet_1_0__leaf_net287),
    .S1(net984),
    .X(net297));
 sky130_fd_sc_hd__buf_1 c323 (.A(clknet_1_0__leaf_net814),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(clknet_1_0__leaf_net298),
    .A1(clknet_1_1__leaf_net273),
    .A2(net288),
    .A3(clknet_1_0__leaf_net287),
    .S0(net286),
    .S1(net147),
    .X(net299));
 sky130_fd_sc_hd__mux4_2 c325 (.A0(clknet_1_1__leaf_net296),
    .A1(net277),
    .A2(net168),
    .A3(net288),
    .S0(net989),
    .S1(net157),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net295),
    .A1(clknet_1_1__leaf_net298),
    .A2(clknet_1_0__leaf_net300),
    .A3(net284),
    .S0(clknet_1_0__leaf_net287),
    .S1(net1004),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(clknet_1_0__leaf_net300),
    .A1(clknet_1_1__leaf_net287),
    .A2(clknet_1_0__leaf_net290),
    .A3(clknet_1_0__leaf_net814),
    .S0(net839),
    .S1(net840),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(clknet_1_0__leaf_net300),
    .A1(clknet_1_0__leaf_net296),
    .A2(clknet_1_1__leaf_net287),
    .A3(net1002),
    .S0(net840),
    .S1(net841),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 c329 (.A0(net303),
    .A1(clknet_1_1__leaf_net287),
    .A2(net269),
    .A3(net266),
    .S0(net840),
    .S1(net841),
    .X(net304));
 sky130_fd_sc_hd__buf_4 c33 (.A(net940),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 c330 (.A(net741),
    .X(net305));
 sky130_fd_sc_hd__xnor2_4 c331 (.A(net305),
    .B(net24),
    .Y(net306));
 sky130_fd_sc_hd__xnor2_1 c332 (.A(net54),
    .B(net841),
    .Y(net307));
 sky130_fd_sc_hd__clkbuf_1 c333 (.A(net740),
    .X(net308));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(clknet_1_1__leaf_net287),
    .A2(net284),
    .B1_N(net179),
    .X(net309));
 sky130_fd_sc_hd__xnor2_1 c335 (.A(net269),
    .B(net46),
    .Y(net310));
 sky130_fd_sc_hd__clkbuf_2 c336 (.A(net765),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net267),
    .A1(net306),
    .A2(net284),
    .A3(net177),
    .S0(net937),
    .S1(net984),
    .X(net312));
 sky130_fd_sc_hd__xnor2_1 c338 (.A(net292),
    .B(clknet_1_1__leaf_net287),
    .Y(net313));
 sky130_fd_sc_hd__mux4_2 c339 (.A0(net188),
    .A1(clknet_1_1__leaf_net300),
    .A2(clknet_1_1__leaf_net309),
    .A3(net984),
    .S0(net33),
    .S1(net311),
    .X(net314));
 sky130_fd_sc_hd__a21bo_1 c34 (.A1(net931),
    .A2(net7),
    .B1_N(net0),
    .X(net9));
 sky130_fd_sc_hd__xnor2_1 c340 (.A(clknet_1_1__leaf_net300),
    .B(net311),
    .Y(net315));
 sky130_fd_sc_hd__a41o_1 c341 (.A1(net189),
    .A2(clknet_1_0__leaf_net313),
    .A3(clknet_1_1__leaf_net314),
    .A4(net178),
    .B1(net292),
    .X(net316));
 sky130_fd_sc_hd__mux4_2 c342 (.A0(net179),
    .A1(net33),
    .A2(net311),
    .A3(net190),
    .S0(net177),
    .S1(net305),
    .X(net317));
 sky130_fd_sc_hd__buf_1 c343 (.A(net761),
    .X(net318));
 sky130_fd_sc_hd__xnor2_2 c344 (.A(net318),
    .B(net317),
    .Y(net319));
 sky130_fd_sc_hd__clkbuf_2 c345 (.A(net909),
    .X(net320));
 sky130_fd_sc_hd__xnor2_1 c346 (.A(net312),
    .B(net177),
    .Y(net321));
 sky130_fd_sc_hd__clkbuf_1 c347 (.A(net761),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net322),
    .A1(clknet_1_0__leaf_net315),
    .A2(net321),
    .A3(net190),
    .S0(net306),
    .S1(net310),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net310),
    .A1(net317),
    .A2(net321),
    .A3(net282),
    .S0(clknet_1_1__leaf_net314),
    .S1(net843),
    .X(net324));
 sky130_fd_sc_hd__xnor2_4 c35 (.A(net5),
    .B(net929),
    .Y(net10));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net169),
    .A1(net190),
    .A2(net308),
    .A3(net321),
    .S0(net841),
    .S1(net843),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net258),
    .A1(net179),
    .A2(net190),
    .A3(net807),
    .S0(net842),
    .S1(net845),
    .X(net326));
 sky130_fd_sc_hd__a21bo_1 c352 (.A1(net78),
    .A2(net326),
    .B1_N(net75),
    .X(net327));
 sky130_fd_sc_hd__a31o_1 c353 (.A1(net317),
    .A2(net320),
    .A3(net30),
    .B1(net832),
    .X(net328));
 sky130_fd_sc_hd__a41o_1 c354 (.A1(net284),
    .A2(net306),
    .A3(net163),
    .A4(clknet_1_0__leaf_net313),
    .B1(net971),
    .X(net329));
 sky130_fd_sc_hd__a31o_2 c355 (.A1(net326),
    .A2(net177),
    .A3(net245),
    .B1(net839),
    .X(net330));
 sky130_fd_sc_hd__a41o_1 c356 (.A1(net70),
    .A2(net937),
    .A3(net180),
    .A4(net787),
    .B1(net1004),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 c357 (.A(net902),
    .X(net332));
 sky130_fd_sc_hd__a41o_1 c358 (.A1(net163),
    .A2(net180),
    .A3(net195),
    .A4(clknet_1_1__leaf_net304),
    .B1(net990),
    .X(net333));
 sky130_fd_sc_hd__a41o_1 c359 (.A1(net195),
    .A2(net1006),
    .A3(net54),
    .A4(net332),
    .B1(net327),
    .X(net334));
 sky130_fd_sc_hd__a21bo_1 c36 (.A1(net7),
    .A2(net0),
    .B1_N(net935),
    .X(net11));
 sky130_fd_sc_hd__a31o_1 c360 (.A1(net168),
    .A2(net75),
    .A3(net940),
    .B1(net832),
    .X(net335));
 sky130_fd_sc_hd__a41o_4 c361 (.A1(net152),
    .A2(net332),
    .A3(net993),
    .A4(net984),
    .B1(net834),
    .X(net336));
 sky130_fd_sc_hd__a41o_1 c362 (.A1(net191),
    .A2(net152),
    .A3(net327),
    .A4(net336),
    .B1(net993),
    .X(net337));
 sky130_fd_sc_hd__sdfrtp_2 c363 (.CLK(clknet_4_14_0_clk),
    .D(net332),
    .RESET_B(net1051),
    .SCD(net336),
    .SCE(net993),
    .Q(net338));
 sky130_fd_sc_hd__sdfbbn_1 c364 (.CLK_N(clknet_4_9_0_clk),
    .D(net329),
    .RESET_B(net993),
    .SCD(net330),
    .SCE(net195),
    .SET_B(net1054),
    .Q(net339));
 sky130_fd_sc_hd__sdfbbp_1 c365 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net313),
    .RESET_B(net241),
    .SCD(clknet_1_0__leaf_net333),
    .SCE(net1074),
    .SET_B(clknet_1_1__leaf_net304),
    .Q(net341),
    .Q_N(net340));
 sky130_fd_sc_hd__sdfbbn_2 c366 (.CLK_N(clknet_4_12_0_clk),
    .D(net327),
    .RESET_B(net338),
    .SCD(net317),
    .SCE(net336),
    .SET_B(net993),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(clknet_1_0__leaf_net333),
    .A1(net266),
    .A2(net340),
    .A3(net993),
    .S0(net46),
    .S1(net332),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c368 (.A0(net341),
    .A1(net948),
    .A2(net54),
    .A3(net335),
    .S0(net342),
    .S1(net846),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_1 c369 (.CLK_N(clknet_4_12_0_clk),
    .D(net177),
    .RESET_B(net338),
    .SCD(clknet_1_1__leaf_net314),
    .SCE(net343),
    .SET_B(net13),
    .Q(net347),
    .Q_N(net346));
 sky130_fd_sc_hd__a41o_4 c37 (.A1(net936),
    .A2(net4),
    .A3(net6),
    .A4(net7),
    .B1(net2),
    .X(net12));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net75),
    .A1(net948),
    .A2(net347),
    .A3(net180),
    .S0(net284),
    .S1(net208),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(net348),
    .A1(net338),
    .A2(net330),
    .A3(net346),
    .S0(net805),
    .S1(net831),
    .X(net349));
 sky130_fd_sc_hd__sdfbbp_1 c372 (.CLK(clknet_4_9_0_clk),
    .D(net347),
    .RESET_B(net336),
    .SCD(net328),
    .SCE(net1059),
    .SET_B(net1050),
    .Q(net350));
 sky130_fd_sc_hd__sdfbbn_1 c373 (.CLK_N(clknet_4_9_0_clk),
    .D(net331),
    .RESET_B(net350),
    .SCD(net948),
    .SCE(clknet_1_1__leaf_net333),
    .SET_B(net1061),
    .Q(net351));
 sky130_fd_sc_hd__a41o_1 c374 (.A1(net223),
    .A2(net229),
    .A3(net209),
    .A4(clknet_1_1__leaf_net290),
    .B1(net950),
    .X(net352));
 sky130_fd_sc_hd__a31o_4 c375 (.A1(net158),
    .A2(net238),
    .A3(net221),
    .B1(net838),
    .X(net353));
 sky130_fd_sc_hd__sdfbbn_1 c376 (.CLK_N(clknet_4_14_0_clk),
    .D(net99),
    .RESET_B(net1056),
    .SCD(net353),
    .SCE(clknet_1_0__leaf_net218),
    .SET_B(net967),
    .Q(net355),
    .Q_N(net354));
 sky130_fd_sc_hd__a41o_1 c377 (.A1(clknet_1_0__leaf_net217),
    .A2(net99),
    .A3(net229),
    .A4(net937),
    .B1(net981),
    .X(net356));
 sky130_fd_sc_hd__sdfbbp_1 c378 (.CLK(clknet_4_14_0_clk),
    .D(net158),
    .RESET_B(clknet_1_0__leaf_net217),
    .SCD(net353),
    .SCE(net342),
    .SET_B(clknet_1_0__leaf_net828),
    .Q(net956),
    .Q_N(net357));
 sky130_fd_sc_hd__a41o_4 c379 (.A1(net168),
    .A2(net1083),
    .A3(net87),
    .A4(net785),
    .B1(net836),
    .X(net953));
 sky130_fd_sc_hd__a21bo_4 c38 (.A1(net10),
    .A2(net929),
    .B1_N(net11),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net158),
    .A1(net353),
    .A2(net208),
    .A3(net224),
    .S0(net784),
    .S1(net805),
    .X(net358));
 sky130_fd_sc_hd__a41o_1 c381 (.A1(net93),
    .A2(net215),
    .A3(net357),
    .A4(net237),
    .B1(clknet_1_0__leaf_net828),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net209),
    .A1(net1044),
    .A2(net99),
    .A3(net953),
    .S0(clknet_1_0__leaf_net828),
    .S1(net835),
    .X(net360));
 sky130_fd_sc_hd__sdfbbn_1 c383 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_0__leaf_net218),
    .RESET_B(net1066),
    .SCD(net953),
    .SCE(net342),
    .SET_B(net1053),
    .Q(net361));
 sky130_fd_sc_hd__sdfbbn_1 c384 (.CLK_N(clknet_4_14_0_clk),
    .D(net359),
    .RESET_B(net1045),
    .SCD(net93),
    .SCE(net338),
    .SET_B(net953),
    .Q(net362));
 sky130_fd_sc_hd__a41o_1 c385 (.A1(net355),
    .A2(net231),
    .A3(net353),
    .A4(clknet_1_1__leaf_net315),
    .B1(net98),
    .X(net363));
 sky130_fd_sc_hd__sdfbbp_1 c386 (.CLK(clknet_4_15_0_clk),
    .D(net238),
    .RESET_B(net953),
    .SCD(net209),
    .SCE(net168),
    .SET_B(net1048),
    .Q(net364));
 sky130_fd_sc_hd__sdfbbn_1 c387 (.CLK_N(clknet_4_14_0_clk),
    .D(net345),
    .RESET_B(net953),
    .SCD(net330),
    .SCE(net306),
    .SET_B(net1075),
    .Q(net366),
    .Q_N(net365));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(net364),
    .A1(net361),
    .A2(clknet_1_1__leaf_net218),
    .A3(net953),
    .S0(net353),
    .S1(net93),
    .X(net367));
 sky130_fd_sc_hd__a41o_1 c389 (.A1(net366),
    .A2(net354),
    .A3(net1042),
    .A4(net353),
    .B1(net849),
    .X(net368));
 sky130_fd_sc_hd__a21bo_4 c39 (.A1(net12),
    .A2(net11),
    .B1_N(net9),
    .X(net14));
 sky130_fd_sc_hd__a31o_1 c390 (.A1(net1042),
    .A2(net209),
    .A3(net957),
    .B1(net353),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net330),
    .A1(net54),
    .A2(clknet_1_1__leaf_net368),
    .A3(net981),
    .S0(net365),
    .S1(net836),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net87),
    .A1(net362),
    .A2(net365),
    .A3(net168),
    .S0(clknet_1_1__leaf_net368),
    .S1(net953),
    .X(net371));
 sky130_fd_sc_hd__sdfbbn_1 c393 (.CLK_N(clknet_4_14_0_clk),
    .D(net338),
    .RESET_B(net366),
    .SCD(net306),
    .SCE(net330),
    .SET_B(clknet_1_1__leaf_net850),
    .Q(net372));
 sky130_fd_sc_hd__a41o_1 c394 (.A1(net369),
    .A2(net366),
    .A3(clknet_1_1__leaf_net368),
    .A4(clknet_1_1__leaf_net850),
    .B1(clknet_1_0__leaf_net851),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net229),
    .A1(net373),
    .A2(net87),
    .A3(clknet_1_1__leaf_net218),
    .S0(net981),
    .S1(clknet_1_1__leaf_net851),
    .X(net374));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net934),
    .B(net241),
    .Y(net375));
 sky130_fd_sc_hd__a21bo_2 c397 (.A1(net126),
    .A2(net259),
    .B1_N(net110),
    .X(net376));
 sky130_fd_sc_hd__xnor2_1 c398 (.A(net1008),
    .B(net375),
    .Y(net377));
 sky130_fd_sc_hd__xnor2_2 c399 (.A(net1001),
    .B(net376),
    .Y(net378));
 sky130_fd_sc_hd__a41o_4 c40 (.A1(net937),
    .A2(net7),
    .A3(net3),
    .A4(net14),
    .B1(net668),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 c400 (.A(net751),
    .X(net379));
 sky130_fd_sc_hd__xnor2_4 c401 (.A(net1000),
    .B(net979),
    .Y(net380));
 sky130_fd_sc_hd__xnor2_1 c402 (.A(net942),
    .B(net248),
    .Y(net381));
 sky130_fd_sc_hd__xnor2_4 c403 (.A(net927),
    .B(net375),
    .Y(net382));
 sky130_fd_sc_hd__clkbuf_4 c404 (.A(net751),
    .X(net383));
 sky130_fd_sc_hd__a21bo_2 c405 (.A1(net379),
    .A2(net375),
    .B1_N(net383),
    .X(net384));
 sky130_fd_sc_hd__xnor2_2 c406 (.A(net377),
    .B(net382),
    .Y(net385));
 sky130_fd_sc_hd__xnor2_4 c407 (.A(net248),
    .B(net380),
    .Y(net386));
 sky130_fd_sc_hd__a21bo_1 c408 (.A1(net110),
    .A2(net1001),
    .B1_N(net375),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 c409 (.A(net1071),
    .X(net388));
 sky130_fd_sc_hd__xnor2_2 c41 (.A(net939),
    .B(net14),
    .Y(net16));
 sky130_fd_sc_hd__a41o_2 c410 (.A1(net384),
    .A2(net386),
    .A3(net108),
    .A4(net382),
    .B1(net971),
    .X(net389));
 sky130_fd_sc_hd__a31o_4 c411 (.A1(net382),
    .A2(net241),
    .A3(net375),
    .B1(net383),
    .X(net390));
 sky130_fd_sc_hd__a21bo_1 c412 (.A1(net381),
    .A2(net383),
    .B1_N(net382),
    .X(net391));
 sky130_fd_sc_hd__a31o_1 c413 (.A1(net386),
    .A2(net389),
    .A3(net384),
    .B1(net391),
    .X(net392));
 sky130_fd_sc_hd__a21bo_1 c414 (.A1(net382),
    .A2(net383),
    .B1_N(net818),
    .X(net393));
 sky130_fd_sc_hd__a31o_1 c415 (.A1(net375),
    .A2(net391),
    .A3(net393),
    .B1(net390),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net388),
    .A1(net384),
    .A2(net247),
    .A3(net389),
    .S0(net382),
    .S1(net391),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net113),
    .A1(net394),
    .A2(net108),
    .A3(net386),
    .S0(net382),
    .S1(net818),
    .X(net396));
 sky130_fd_sc_hd__xnor2_2 c418 (.A(net390),
    .B(net255),
    .Y(net397));
 sky130_fd_sc_hd__xnor2_2 c419 (.A(net134),
    .B(net983),
    .Y(net398));
 sky130_fd_sc_hd__a41o_1 c42 (.A1(net16),
    .A2(net14),
    .A3(net11),
    .A4(net9),
    .B1(net2),
    .X(net17));
 sky130_fd_sc_hd__xnor2_2 c420 (.A(net247),
    .B(net384),
    .Y(net399));
 sky130_fd_sc_hd__xnor2_2 c421 (.A(net1001),
    .B(net387),
    .Y(net400));
 sky130_fd_sc_hd__xnor2_2 c422 (.A(net271),
    .B(net817),
    .Y(net401));
 sky130_fd_sc_hd__xnor2_4 c423 (.A(net994),
    .B(net818),
    .Y(net402));
 sky130_fd_sc_hd__xnor2_1 c424 (.A(net258),
    .B(net144),
    .Y(net403));
 sky130_fd_sc_hd__a21bo_1 c425 (.A1(net398),
    .A2(net983),
    .B1_N(net400),
    .X(net404));
 sky130_fd_sc_hd__xnor2_1 c426 (.A(net402),
    .B(net404),
    .Y(net405));
 sky130_fd_sc_hd__buf_1 c427 (.A(net796),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net401),
    .A1(net402),
    .A2(net390),
    .A3(net123),
    .S0(net282),
    .S1(net983),
    .X(net407));
 sky130_fd_sc_hd__a41o_1 c429 (.A1(net144),
    .A2(clknet_1_0__leaf_net279),
    .A3(net400),
    .A4(net983),
    .B1(net818),
    .X(net408));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net16),
    .A1(net935),
    .A2(net12),
    .A3(net14),
    .S0(net1),
    .S1(net989),
    .X(net18));
 sky130_fd_sc_hd__xnor2_2 c430 (.A(net261),
    .B(net401),
    .Y(net409));
 sky130_fd_sc_hd__xnor2_1 c431 (.A(net405),
    .B(clknet_1_0__leaf_net408),
    .Y(net964));
 sky130_fd_sc_hd__a21bo_1 c432 (.A1(net403),
    .A2(net387),
    .B1_N(clknet_1_0__leaf_net964),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net145),
    .A1(net404),
    .A2(net965),
    .A3(net398),
    .S0(clknet_1_0__leaf_net964),
    .S1(net951),
    .X(net411));
 sky130_fd_sc_hd__a21bo_1 c434 (.A1(net255),
    .A2(net399),
    .B1_N(clknet_1_0__leaf_net964),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 c435 (.A(net796),
    .X(net413));
 sky130_fd_sc_hd__sdfsbp_1 c436 (.CLK(clknet_4_5_0_clk),
    .D(net278),
    .SCD(clknet_1_0__leaf_net411),
    .SCE(net409),
    .SET_B(clknet_1_0__leaf_net964),
    .Q(net415),
    .Q_N(net414));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_0__leaf_net410),
    .A1(net405),
    .A2(clknet_1_0__leaf_net412),
    .A3(net983),
    .S0(net415),
    .S1(net402),
    .X(net416));
 sky130_fd_sc_hd__sdfsbp_2 c438 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net412),
    .SCD(clknet_1_1__leaf_net410),
    .SCE(net1062),
    .SET_B(clknet_1_0__leaf_net964),
    .Q(net418),
    .Q_N(net417));
 sky130_fd_sc_hd__buf_1 c439 (.A(net796),
    .X(net419));
 sky130_fd_sc_hd__xnor2_4 c44 (.A(net1047),
    .B(net997),
    .Y(net19));
 sky130_fd_sc_hd__sdfbbp_1 c440 (.CLK(clknet_4_4_0_clk),
    .D(net447),
    .RESET_B(net22),
    .SCD(net384),
    .SCE(net970),
    .SET_B(net979),
    .Q(net421),
    .Q_N(net420));
 sky130_fd_sc_hd__buf_2 c441 (.A(net900),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 c442 (.A(net900),
    .X(net423));
 sky130_fd_sc_hd__sdfbbn_2 c443 (.CLK_N(clknet_4_4_0_clk),
    .D(net422),
    .RESET_B(net389),
    .SCD(net420),
    .SCE(clknet_1_0__leaf_net304),
    .SET_B(clknet_1_0__leaf_net964),
    .Q(net425),
    .Q_N(net424));
 sky130_fd_sc_hd__a41o_1 c444 (.A1(net399),
    .A2(net425),
    .A3(net133),
    .A4(net422),
    .B1(net241),
    .X(net426));
 sky130_fd_sc_hd__sdfbbn_1 c445 (.CLK_N(clknet_4_6_0_clk),
    .D(net421),
    .RESET_B(net423),
    .SCD(net258),
    .SCE(net422),
    .SET_B(clknet_1_0__leaf_net290),
    .Q(net428),
    .Q_N(net427));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net262),
    .A1(net446),
    .A2(net422),
    .A3(net421),
    .S0(net970),
    .S1(net854),
    .X(net429));
 sky130_fd_sc_hd__sdfbbp_1 c447 (.CLK(clknet_4_4_0_clk),
    .D(net441),
    .RESET_B(net445),
    .SCD(net406),
    .SCE(net425),
    .SET_B(net1057),
    .Q(net431),
    .Q_N(net430));
 sky130_fd_sc_hd__sdfbbn_1 c448 (.CLK_N(clknet_4_4_0_clk),
    .D(net22),
    .RESET_B(net970),
    .SCD(net422),
    .SCE(net430),
    .SET_B(net857),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net150),
    .A1(net419),
    .A2(net285),
    .A3(net1002),
    .S0(net422),
    .S1(net430),
    .X(net434));
 sky130_fd_sc_hd__xnor2_4 c45 (.A(net989),
    .B(net40),
    .Y(net20));
 sky130_fd_sc_hd__a41o_1 c450 (.A1(net990),
    .A2(net418),
    .A3(clknet_1_0__leaf_net304),
    .A4(net970),
    .B1(net817),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(net431),
    .A1(net422),
    .A2(net432),
    .A3(net419),
    .S0(clknet_1_1__leaf_net964),
    .S1(clknet_1_0__leaf_net816),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(clknet_1_0__leaf_net273),
    .A1(net421),
    .A2(net970),
    .A3(net983),
    .S0(net787),
    .S1(net855),
    .X(net437));
 sky130_fd_sc_hd__a41o_1 c453 (.A1(clknet_1_0__leaf_net436),
    .A2(net159),
    .A3(net422),
    .A4(net18),
    .B1(net856),
    .X(net438));
 sky130_fd_sc_hd__a21bo_1 c454 (.A1(net406),
    .A2(net431),
    .B1_N(net428),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net998),
    .A1(clknet_1_1__leaf_net436),
    .A2(net282),
    .A3(net1002),
    .S0(net430),
    .S1(clknet_1_1__leaf_net816),
    .X(net440));
 sky130_fd_sc_hd__a21bo_1 c456 (.A1(clknet_1_1__leaf_net279),
    .A2(clknet_1_0__leaf_net408),
    .B1_N(net266),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net137),
    .A1(net409),
    .A2(net406),
    .A3(net285),
    .S0(clknet_1_0__leaf_net304),
    .S1(net417),
    .X(net442));
 sky130_fd_sc_hd__a21bo_1 c458 (.A1(net930),
    .A2(net266),
    .B1_N(net22),
    .X(net443));
 sky130_fd_sc_hd__a41o_1 c459 (.A1(clknet_1_0__leaf_net304),
    .A2(net990),
    .A3(clknet_1_0__leaf_net964),
    .A4(net817),
    .B1(net855),
    .X(net444));
 sky130_fd_sc_hd__xnor2_4 c46 (.A(net668),
    .B(net923),
    .Y(net21));
 sky130_fd_sc_hd__a21bo_1 c460 (.A1(net133),
    .A2(net285),
    .B1_N(net282),
    .X(net445));
 sky130_fd_sc_hd__sdfbbn_1 c461 (.CLK_N(clknet_4_4_0_clk),
    .D(net404),
    .RESET_B(net262),
    .SCD(net418),
    .SCE(net970),
    .SET_B(net983),
    .Q(net447),
    .Q_N(net446));
 sky130_fd_sc_hd__a21bo_4 c462 (.A1(net413),
    .A2(net443),
    .B1_N(net984),
    .X(net448));
 sky130_fd_sc_hd__a21bo_1 c463 (.A1(net431),
    .A2(net998),
    .B1_N(net282),
    .X(net449));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(net925),
    .A1(net258),
    .A2(net186),
    .A3(net423),
    .S0(net448),
    .S1(net965),
    .X(net450));
 sky130_fd_sc_hd__a31o_1 c465 (.A1(net449),
    .A2(net24),
    .A3(net320),
    .B1(net430),
    .X(net451));
 sky130_fd_sc_hd__sdfstp_1 c466 (.CLK(clknet_4_9_0_clk),
    .D(net311),
    .SCD(net451),
    .SCE(net320),
    .SET_B(net990),
    .Q(net960));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_0__leaf_net290),
    .A1(net282),
    .A2(net431),
    .A3(net1002),
    .S0(net319),
    .S1(net818),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net57),
    .A1(net311),
    .A2(clknet_1_1__leaf_net964),
    .A3(clknet_1_0__leaf_net290),
    .S0(net842),
    .S1(net859),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net282),
    .A1(net319),
    .A2(clknet_1_1__leaf_net314),
    .A3(clknet_1_1__leaf_net408),
    .S0(net817),
    .S1(net861),
    .X(net454));
 sky130_fd_sc_hd__a21bo_4 c47 (.A1(net9),
    .A2(net20),
    .B1_N(net942),
    .X(net22));
 sky130_fd_sc_hd__sdfstp_2 c470 (.CLK(clknet_4_9_0_clk),
    .D(net451),
    .SCD(net311),
    .SCE(clknet_1_0__leaf_net315),
    .SET_B(net860),
    .Q(net455));
 sky130_fd_sc_hd__a41o_1 c471 (.A1(clknet_1_0__leaf_net304),
    .A2(net455),
    .A3(net24),
    .A4(net802),
    .B1(net860),
    .X(net456));
 sky130_fd_sc_hd__buf_1 c472 (.A(net899),
    .X(net457));
 sky130_fd_sc_hd__a21bo_1 c473 (.A1(clknet_1_0__leaf_net408),
    .A2(net1002),
    .B1_N(net457),
    .X(net458));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(clknet_1_1__leaf_net456),
    .A2(net245),
    .B1_N(net990),
    .X(net459));
 sky130_fd_sc_hd__a41o_1 c475 (.A1(clknet_1_1__leaf_net459),
    .A2(net960),
    .A3(clknet_1_1__leaf_net964),
    .A4(net842),
    .B1(net845),
    .X(net460));
 sky130_fd_sc_hd__a21bo_1 c476 (.A1(net457),
    .A2(net431),
    .B1_N(net269),
    .X(net461));
 sky130_fd_sc_hd__a21bo_1 c477 (.A1(net285),
    .A2(net428),
    .B1_N(clknet_1_0__leaf_net459),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net458),
    .A1(clknet_1_0__leaf_net462),
    .A2(net178),
    .A3(net970),
    .S0(net450),
    .S1(net397),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net245),
    .A1(net455),
    .A2(clknet_1_0__leaf_net459),
    .A3(net449),
    .S0(net802),
    .S1(net861),
    .X(net464));
 sky130_fd_sc_hd__xnor2_4 c48 (.A(net1018),
    .B(net21),
    .Y(net23));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(clknet_1_1__leaf_net464),
    .A1(net461),
    .A2(clknet_1_0__leaf_net456),
    .A3(clknet_1_0__leaf_net290),
    .S0(clknet_1_1__leaf_net964),
    .S1(net801),
    .X(net465));
 sky130_fd_sc_hd__buf_1 c481 (.A(net898),
    .X(net466));
 sky130_fd_sc_hd__a21bo_1 c482 (.A1(net843),
    .A2(net861),
    .B1_N(net863),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net57),
    .A1(net457),
    .A2(net467),
    .A3(net970),
    .S0(net461),
    .S1(clknet_1_1__leaf_net964),
    .X(net468));
 sky130_fd_sc_hd__xnor2_1 c484 (.A(net926),
    .B(net343),
    .Y(net469));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net328),
    .A1(net455),
    .A2(net423),
    .A3(clknet_1_1__leaf_net304),
    .S0(net186),
    .S1(net990),
    .X(net470));
 sky130_fd_sc_hd__xnor2_1 c486 (.A(net944),
    .B(net466),
    .Y(net471));
 sky130_fd_sc_hd__a21bo_2 c487 (.A1(net423),
    .A2(net306),
    .B1_N(net846),
    .X(net472));
 sky130_fd_sc_hd__xnor2_1 c488 (.A(clknet_1_1__leaf_net304),
    .B(net472),
    .Y(net473));
 sky130_fd_sc_hd__a31o_1 c489 (.A1(net450),
    .A2(net1006),
    .A3(net980),
    .B1(net245),
    .X(net474));
 sky130_fd_sc_hd__xnor2_4 c49 (.A(net1029),
    .B(net936),
    .Y(net24));
 sky130_fd_sc_hd__xnor2_1 c490 (.A(net423),
    .B(net245),
    .Y(net475));
 sky130_fd_sc_hd__xnor2_1 c491 (.A(net971),
    .B(net862),
    .Y(net476));
 sky130_fd_sc_hd__a21bo_1 c492 (.A1(net992),
    .A2(net46),
    .B1_N(net948),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net339),
    .A1(net450),
    .A2(net472),
    .A3(clknet_1_1__leaf_net304),
    .S0(net336),
    .S1(net823),
    .X(net478));
 sky130_fd_sc_hd__a21bo_1 c494 (.A1(net993),
    .A2(net820),
    .B1_N(net866),
    .X(net479));
 sky130_fd_sc_hd__a21bo_1 c495 (.A1(net474),
    .A2(clknet_1_0__leaf_net315),
    .B1_N(net841),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 c496 (.A(net750),
    .X(net481));
 sky130_fd_sc_hd__buf_1 c497 (.A(net902),
    .X(net949));
 sky130_fd_sc_hd__buf_1 c498 (.A(net750),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 c499 (.A(net759),
    .X(net483));
 sky130_fd_sc_hd__xnor2_2 c50 (.A(net927),
    .B(net22),
    .Y(net25));
 sky130_fd_sc_hd__clkbuf_1 c500 (.A(net760),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net384),
    .A1(net483),
    .A2(net328),
    .A3(clknet_1_0__leaf_net315),
    .S0(net482),
    .S1(net866),
    .X(net485));
 sky130_fd_sc_hd__a21bo_1 c502 (.A1(net320),
    .A2(net481),
    .B1_N(clknet_1_1__leaf_net473),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net486),
    .A1(net993),
    .A2(net482),
    .A3(clknet_1_1__leaf_net304),
    .S0(net336),
    .S1(net867),
    .X(net487));
 sky130_fd_sc_hd__buf_1 c504 (.A(clknet_1_1__leaf_net903),
    .X(net488));
 sky130_fd_sc_hd__a21bo_1 c505 (.A1(net488),
    .A2(net474),
    .B1_N(net819),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c509 (.A0(clknet_1_1__leaf_net290),
    .A1(net472),
    .A2(net981),
    .A3(net427),
    .S0(net950),
    .S1(net852),
    .X(net490));
 sky130_fd_sc_hd__xnor2_4 c51 (.A(net1028),
    .B(net3),
    .Y(net26));
 sky130_fd_sc_hd__mux4_1 c510 (.A0(net30),
    .A1(net19),
    .A2(net1032),
    .A3(net472),
    .S0(net950),
    .S1(clknet_1_0__leaf_net850),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c511 (.A0(net981),
    .A1(net967),
    .A2(net966),
    .A3(net472),
    .S0(net214),
    .S1(net952),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c512 (.A0(net1005),
    .A1(net353),
    .A2(net960),
    .A3(clknet_1_1__leaf_net290),
    .S0(net957),
    .S1(clknet_1_0__leaf_net368),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c513 (.A0(net306),
    .A1(clknet_1_1__leaf_net408),
    .A2(clknet_1_1__leaf_net290),
    .A3(net981),
    .S0(net958),
    .S1(net357),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c514 (.A0(clknet_1_1__leaf_net368),
    .A1(clknet_1_1__leaf_net491),
    .A2(net956),
    .A3(net967),
    .S0(net981),
    .S1(clknet_1_1__leaf_net315),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c515 (.A0(net372),
    .A1(net1019),
    .A2(clknet_1_1__leaf_net315),
    .A3(net342),
    .S0(net953),
    .S1(clknet_1_1__leaf_net850),
    .X(net496));
 sky130_fd_sc_hd__mux4_2 c516 (.A0(net937),
    .A1(net967),
    .A2(net343),
    .A3(net214),
    .S0(net789),
    .S1(net853),
    .X(net969));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(clknet_1_1__leaf_net315),
    .A1(net971),
    .A2(net342),
    .A3(net822),
    .S0(net863),
    .S1(clknet_1_0__leaf_net869),
    .X(net497));
 sky130_fd_sc_hd__mux4_2 c518 (.A0(net472),
    .A1(net363),
    .A2(net306),
    .A3(net427),
    .S0(net353),
    .S1(net955),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(clknet_1_1__leaf_net498),
    .A1(net343),
    .A2(net981),
    .A3(clknet_1_0__leaf_net850),
    .S0(net868),
    .S1(clknet_1_1__leaf_net869),
    .X(net499));
 sky130_fd_sc_hd__xnor2_4 c52 (.A(net982),
    .B(net942),
    .Y(net27));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(net358),
    .A1(net953),
    .A2(net922),
    .A3(clknet_1_0__leaf_net368),
    .S0(clknet_1_1__leaf_net499),
    .S1(clknet_1_0__leaf_net963),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(net232),
    .A1(net492),
    .A2(clknet_1_0__leaf_net491),
    .A3(clknet_1_1__leaf_net499),
    .S0(clknet_1_1__leaf_net290),
    .S1(clknet_1_0__leaf_net963),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net475),
    .A1(clknet_1_1__leaf_net964),
    .A2(clknet_1_0__leaf_net499),
    .A3(net1005),
    .S0(clknet_1_0__leaf_net368),
    .S1(net861),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net343),
    .A1(net497),
    .A2(net967),
    .A3(clknet_1_1__leaf_net499),
    .S0(net260),
    .S1(net955),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(clknet_1_1__leaf_net502),
    .A1(net1005),
    .A2(net948),
    .A3(net472),
    .S0(net870),
    .S1(net872),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(clknet_1_0__leaf_net498),
    .A1(clknet_1_0__leaf_net499),
    .A2(net467),
    .A3(clknet_1_0__leaf_net368),
    .S0(net950),
    .S1(clknet_1_0__leaf_net869),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net467),
    .A1(clknet_1_0__leaf_net502),
    .A2(net343),
    .A3(clknet_1_1__leaf_net315),
    .S0(net984),
    .S1(net871),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net23),
    .A1(net428),
    .A2(net505),
    .A3(net969),
    .S0(clknet_1_0__leaf_net491),
    .S1(clknet_1_0__leaf_net499),
    .X(net507));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net987),
    .B(net976),
    .Y(net508));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net383),
    .B(net976),
    .Y(net509));
 sky130_fd_sc_hd__xnor2_4 c53 (.A(net934),
    .B(net997),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_1 c530 (.A(net971),
    .B(net1000),
    .Y(net510));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net385),
    .B(net1000),
    .Y(net511));
 sky130_fd_sc_hd__clkbuf_1 c532 (.A(net729),
    .X(net512));
 sky130_fd_sc_hd__xnor2_1 c533 (.A(net383),
    .B(net508),
    .Y(net513));
 sky130_fd_sc_hd__buf_1 c534 (.A(net729),
    .X(net514));
 sky130_fd_sc_hd__xnor2_4 c535 (.A(net509),
    .B(net508),
    .Y(net515));
 sky130_fd_sc_hd__xnor2_1 c536 (.A(net959),
    .B(net971),
    .Y(net516));
 sky130_fd_sc_hd__dlymetal6s2s_1 c537 (.A(net800),
    .X(net517));
 sky130_fd_sc_hd__buf_4 c538 (.A(net800),
    .X(net518));
 sky130_fd_sc_hd__buf_1 c539 (.A(net912),
    .X(net519));
 sky130_fd_sc_hd__xnor2_4 c54 (.A(net943),
    .B(net26),
    .Y(net29));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(net396),
    .A2(net519),
    .B1_N(net509),
    .X(net520));
 sky130_fd_sc_hd__xnor2_1 c541 (.A(net938),
    .B(net511),
    .Y(net521));
 sky130_fd_sc_hd__clkbuf_1 c542 (.A(net912),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 c543 (.A(net799),
    .X(net523));
 sky130_fd_sc_hd__xnor2_1 c544 (.A(net522),
    .B(net517),
    .Y(net524));
 sky130_fd_sc_hd__a21bo_1 c545 (.A1(net514),
    .A2(net519),
    .B1_N(net511),
    .X(net525));
 sky130_fd_sc_hd__xnor2_2 c546 (.A(net524),
    .B(net514),
    .Y(net526));
 sky130_fd_sc_hd__a31o_1 c547 (.A1(net519),
    .A2(net523),
    .A3(net526),
    .B1(net509),
    .X(net527));
 sky130_fd_sc_hd__a21bo_4 c548 (.A1(net527),
    .A2(net525),
    .B1_N(net517),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net517),
    .A1(net527),
    .A2(net526),
    .A3(net528),
    .S0(net523),
    .S1(net512),
    .X(net529));
 sky130_fd_sc_hd__mux4_2 c55 (.A0(net23),
    .A1(net2),
    .A2(net9),
    .A3(net18),
    .S0(net29),
    .S1(net997),
    .X(net30));
 sky130_fd_sc_hd__xnor2_1 c550 (.A(net994),
    .B(net523),
    .Y(net530));
 sky130_fd_sc_hd__a21bo_2 c551 (.A1(net509),
    .A2(net387),
    .B1_N(net518),
    .X(net531));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net937),
    .A1(net525),
    .A2(net994),
    .A3(net509),
    .S0(net18),
    .S1(clknet_1_0__leaf_net964),
    .X(net532));
 sky130_fd_sc_hd__xnor2_1 c553 (.A(net18),
    .B(net376),
    .Y(net533));
 sky130_fd_sc_hd__a21bo_1 c554 (.A1(net10),
    .A2(net402),
    .B1_N(net123),
    .X(net534));
 sky130_fd_sc_hd__xnor2_1 c555 (.A(net530),
    .B(net241),
    .Y(net535));
 sky130_fd_sc_hd__a21bo_1 c556 (.A1(net142),
    .A2(net390),
    .B1_N(net531),
    .X(net536));
 sky130_fd_sc_hd__buf_2 c557 (.A(net735),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net523),
    .A1(net515),
    .A2(net415),
    .A3(net979),
    .S0(net397),
    .S1(net534),
    .X(net538));
 sky130_fd_sc_hd__buf_2 c559 (.A(net735),
    .X(net539));
 sky130_fd_sc_hd__a21bo_2 c56 (.A1(net28),
    .A2(net40),
    .B1_N(net29),
    .X(net31));
 sky130_fd_sc_hd__buf_1 c560 (.A(net799),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 c561 (.A(net806),
    .X(net541));
 sky130_fd_sc_hd__buf_1 c562 (.A(net916),
    .X(net542));
 sky130_fd_sc_hd__mux4_2 c563 (.A0(net387),
    .A1(net540),
    .A2(net1000),
    .A3(net415),
    .S0(net537),
    .S1(net541),
    .X(net543));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net538),
    .A1(net542),
    .A2(net274),
    .A3(net540),
    .S0(net537),
    .S1(clknet_1_0__leaf_net964),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 c565 (.A(net779),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net274),
    .A1(net537),
    .A2(net536),
    .A3(net509),
    .S0(net531),
    .S1(net543),
    .X(net546));
 sky130_fd_sc_hd__a31o_4 c567 (.A1(net539),
    .A2(net537),
    .A3(net806),
    .B1(net874),
    .X(net954));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net533),
    .A1(net400),
    .A2(net954),
    .A3(net536),
    .S0(net543),
    .S1(net874),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_2 c569 (.A(net914),
    .X(net548));
 sky130_fd_sc_hd__xnor2_4 c57 (.A(net29),
    .B(net28),
    .Y(net32));
 sky130_fd_sc_hd__a21bo_1 c570 (.A1(net141),
    .A2(net548),
    .B1_N(net875),
    .X(net549));
 sky130_fd_sc_hd__xnor2_1 c571 (.A(net549),
    .B(net875),
    .Y(net550));
 sky130_fd_sc_hd__xnor2_1 c572 (.A(net159),
    .B(net425),
    .Y(net551));
 sky130_fd_sc_hd__clkbuf_1 c573 (.A(net744),
    .X(net552));
 sky130_fd_sc_hd__xnor2_2 c574 (.A(net518),
    .B(net1004),
    .Y(net553));
 sky130_fd_sc_hd__xnor2_1 c575 (.A(net525),
    .B(net439),
    .Y(net554));
 sky130_fd_sc_hd__a31o_2 c576 (.A1(net543),
    .A2(net425),
    .A3(net37),
    .B1(net858),
    .X(net555));
 sky130_fd_sc_hd__a21bo_1 c577 (.A1(net425),
    .A2(net534),
    .B1_N(net873),
    .X(net556));
 sky130_fd_sc_hd__a21bo_2 c578 (.A1(net534),
    .A2(net555),
    .B1_N(net875),
    .X(net557));
 sky130_fd_sc_hd__a41o_1 c579 (.A1(net37),
    .A2(clknet_1_0__leaf_net964),
    .A3(net424),
    .A4(net557),
    .B1(net18),
    .X(net558));
 sky130_fd_sc_hd__a31o_4 c58 (.A1(net1021),
    .A2(net32),
    .A3(net28),
    .B1(net9),
    .X(net33));
 sky130_fd_sc_hd__buf_1 c580 (.A(net743),
    .X(net559));
 sky130_fd_sc_hd__a21bo_1 c581 (.A1(net552),
    .A2(net559),
    .B1_N(net787),
    .X(net560));
 sky130_fd_sc_hd__a21bo_4 c582 (.A1(net560),
    .A2(net130),
    .B1_N(net873),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 c583 (.A(net1049),
    .X(net562));
 sky130_fd_sc_hd__a21bo_1 c584 (.A1(net539),
    .A2(net266),
    .B1_N(net858),
    .X(net563));
 sky130_fd_sc_hd__mux4_2 c585 (.A0(net983),
    .A1(net553),
    .A2(net543),
    .A3(net555),
    .S0(net998),
    .S1(net793),
    .X(net564));
 sky130_fd_sc_hd__a21bo_1 c586 (.A1(net563),
    .A2(net560),
    .B1_N(net561),
    .X(net565));
 sky130_fd_sc_hd__a21bo_2 c587 (.A1(net130),
    .A2(net553),
    .B1_N(net874),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net565),
    .A1(net531),
    .A2(net566),
    .A3(net551),
    .S0(net560),
    .S1(net250),
    .X(net567));
 sky130_fd_sc_hd__sdfbbp_1 c589 (.CLK(clknet_4_3_0_clk),
    .D(net433),
    .RESET_B(net426),
    .SCD(net557),
    .SCE(net30),
    .SET_B(net998),
    .Q(net568));
 sky130_fd_sc_hd__xnor2_2 c59 (.A(net32),
    .B(net1084),
    .Y(net34));
 sky130_fd_sc_hd__a21bo_4 c590 (.A1(net566),
    .A2(net561),
    .B1_N(net792),
    .X(net569));
 sky130_fd_sc_hd__xnor2_4 c591 (.A(net566),
    .B(net569),
    .Y(net570));
 sky130_fd_sc_hd__a41o_1 c592 (.A1(net568),
    .A2(net555),
    .A3(net566),
    .A4(net570),
    .B1(net561),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net562),
    .A1(net561),
    .A2(net570),
    .A3(net424),
    .S0(net551),
    .S1(net922),
    .X(net572));
 sky130_fd_sc_hd__buf_1 c594 (.A(net901),
    .X(net573));
 sky130_fd_sc_hd__a21bo_1 c595 (.A1(net553),
    .A2(net823),
    .B1_N(net862),
    .X(net574));
 sky130_fd_sc_hd__a21bo_1 c596 (.A1(net555),
    .A2(net999),
    .B1_N(net862),
    .X(net575));
 sky130_fd_sc_hd__buf_1 c597 (.A(net901),
    .X(net576));
 sky130_fd_sc_hd__a21bo_1 c598 (.A1(net1002),
    .A2(net965),
    .B1_N(net822),
    .X(net577));
 sky130_fd_sc_hd__a21bo_1 c599 (.A1(net241),
    .A2(net569),
    .B1_N(net576),
    .X(net578));
 sky130_fd_sc_hd__xnor2_4 c60 (.A(net1046),
    .B(net1020),
    .Y(net35));
 sky130_fd_sc_hd__a21bo_1 c600 (.A1(net577),
    .A2(net1077),
    .B1_N(net865),
    .X(net579));
 sky130_fd_sc_hd__buf_1 c601 (.A(clknet_1_0__leaf_net903),
    .X(net580));
 sky130_fd_sc_hd__a21bo_1 c602 (.A1(net999),
    .A2(net1004),
    .B1_N(net865),
    .X(net581));
 sky130_fd_sc_hd__buf_1 c603 (.A(clknet_1_0__leaf_net904),
    .X(net582));
 sky130_fd_sc_hd__sdfbbn_1 c604 (.CLK_N(clknet_4_3_0_clk),
    .D(net389),
    .RESET_B(clknet_1_0__leaf_net580),
    .SCD(clknet_1_0__leaf_net462),
    .SCE(net424),
    .SET_B(net874),
    .Q(net584),
    .Q_N(net583));
 sky130_fd_sc_hd__buf_1 c605 (.A(clknet_1_1__leaf_net904),
    .X(net585));
 sky130_fd_sc_hd__a21bo_1 c606 (.A1(net425),
    .A2(net584),
    .B1_N(clknet_1_0__leaf_net580),
    .X(net586));
 sky130_fd_sc_hd__a21bo_1 c607 (.A1(net585),
    .A2(net555),
    .B1_N(clknet_1_1__leaf_net580),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net574),
    .A1(net561),
    .A2(net999),
    .A3(net571),
    .S0(net448),
    .S1(net874),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_1__leaf_net587),
    .A1(net578),
    .A2(net577),
    .A3(net999),
    .S0(clknet_1_1__leaf_net586),
    .S1(net864),
    .X(net589));
 sky130_fd_sc_hd__xnor2_2 c61 (.A(net932),
    .B(net35),
    .Y(net36));
 sky130_fd_sc_hd__clkbuf_1 c610 (.A(net913),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net542),
    .A1(clknet_1_0__leaf_net586),
    .A2(clknet_1_0__leaf_net580),
    .A3(net999),
    .S0(net980),
    .S1(net424),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net1077),
    .A1(net581),
    .A2(clknet_1_1__leaf_net586),
    .A3(clknet_1_0__leaf_net587),
    .S0(net954),
    .S1(net455),
    .X(net592));
 sky130_fd_sc_hd__a21bo_2 c613 (.A1(net990),
    .A2(net782),
    .B1_N(net876),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_0__leaf_net586),
    .A1(net591),
    .A2(net593),
    .A3(net528),
    .S0(net980),
    .S1(clknet_1_1__leaf_net964),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(clknet_1_1__leaf_net580),
    .A1(net593),
    .A2(clknet_1_1__leaf_net586),
    .A3(net573),
    .S0(net946),
    .S1(net877),
    .X(net595));
 sky130_fd_sc_hd__a31o_1 c616 (.A1(net922),
    .A2(net590),
    .A3(net940),
    .B1(net178),
    .X(net596));
 sky130_fd_sc_hd__sdfbbn_1 c617 (.CLK_N(clknet_4_10_0_clk),
    .D(net186),
    .RESET_B(net479),
    .SCD(net557),
    .SCE(net561),
    .SET_B(net867),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__a31o_1 c618 (.A1(net561),
    .A2(net336),
    .A3(net944),
    .B1(net839),
    .X(net599));
 sky130_fd_sc_hd__a31o_1 c619 (.A1(net448),
    .A2(net993),
    .A3(net455),
    .B1(net180),
    .X(net600));
 sky130_fd_sc_hd__a31o_2 c62 (.A1(net935),
    .A2(net31),
    .A3(net28),
    .B1(net35),
    .X(net37));
 sky130_fd_sc_hd__mux4_2 c620 (.A0(net448),
    .A1(net954),
    .A2(net561),
    .A3(net214),
    .S0(net1004),
    .S1(net862),
    .X(net601));
 sky130_fd_sc_hd__sdfstp_1 c621 (.CLK(clknet_4_10_0_clk),
    .D(net336),
    .SCD(clknet_1_1__leaf_net489),
    .SCE(net482),
    .SET_B(net561),
    .Q(net602));
 sky130_fd_sc_hd__a31o_1 c622 (.A1(net24),
    .A2(net980),
    .A3(net602),
    .B1(net590),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net46),
    .A1(net596),
    .A2(net570),
    .A3(net557),
    .S0(net601),
    .S1(net479),
    .X(net604));
 sky130_fd_sc_hd__a31o_1 c624 (.A1(net1067),
    .A2(net570),
    .A3(net1012),
    .B1(net878),
    .X(net605));
 sky130_fd_sc_hd__a31o_1 c625 (.A1(net993),
    .A2(net215),
    .A3(clknet_1_1__leaf_net964),
    .B1(net808),
    .X(net606));
 sky130_fd_sc_hd__sdfbbp_1 c626 (.CLK(clknet_4_8_0_clk),
    .D(net319),
    .RESET_B(net606),
    .SCD(net477),
    .SCE(net215),
    .SET_B(net879),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__a31o_1 c627 (.A1(net980),
    .A2(net823),
    .A3(net1004),
    .B1(net880),
    .X(net609));
 sky130_fd_sc_hd__sdfbbn_1 c628 (.CLK_N(clknet_4_10_0_clk),
    .D(net482),
    .RESET_B(net605),
    .SCD(net336),
    .SCE(net600),
    .SET_B(net879),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__a31o_4 c629 (.A1(net600),
    .A2(net561),
    .A3(net601),
    .B1(net186),
    .X(net612));
 sky130_fd_sc_hd__a31o_1 c63 (.A1(net2),
    .A2(net34),
    .A3(net35),
    .B1(net37),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net455),
    .A1(net980),
    .A2(net612),
    .A3(net862),
    .S0(net867),
    .S1(net880),
    .X(net613));
 sky130_fd_sc_hd__a41o_1 c631 (.A1(net611),
    .A2(net477),
    .A3(net612),
    .A4(clknet_1_0__leaf_net314),
    .B1(clknet_1_1__leaf_net964),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net1039),
    .A1(net1012),
    .A2(net46),
    .A3(net609),
    .S0(net612),
    .S1(net214),
    .X(net615));
 sky130_fd_sc_hd__sdfbbn_1 c633 (.CLK_N(clknet_4_8_0_clk),
    .D(net180),
    .RESET_B(net557),
    .SCD(net612),
    .SCE(net954),
    .SET_B(net613),
    .Q(net617),
    .Q_N(net616));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net557),
    .A1(clknet_1_0__leaf_net489),
    .A2(net617),
    .A3(net612),
    .S0(net967),
    .S1(net808),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net613),
    .A1(net180),
    .A2(net616),
    .A3(net954),
    .S0(net612),
    .S1(net881),
    .X(net619));
 sky130_fd_sc_hd__mux4_2 c636 (.A0(net615),
    .A1(net617),
    .A2(net180),
    .A3(net612),
    .S0(net1040),
    .S1(net867),
    .X(net945));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net619),
    .A1(net603),
    .A2(net610),
    .A3(net597),
    .S0(net945),
    .S1(net616),
    .X(net620));
 sky130_fd_sc_hd__a41o_1 c64 (.A1(net38),
    .A2(net36),
    .A3(net35),
    .A4(net25),
    .B1(net34),
    .X(net39));
 sky130_fd_sc_hd__xnor2_4 c65 (.A(net2),
    .B(net936),
    .Y(net40));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net31),
    .B(net936),
    .Y(net41));
 sky130_fd_sc_hd__xnor2_1 c660 (.A(net257),
    .B(net390),
    .Y(net621));
 sky130_fd_sc_hd__xnor2_1 c661 (.A(net390),
    .B(net1076),
    .Y(net622));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net386),
    .B(net526),
    .Y(net623));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net393),
    .B(net873),
    .Y(net624));
 sky130_fd_sc_hd__xnor2_4 c664 (.A(net109),
    .B(net518),
    .Y(net625));
 sky130_fd_sc_hd__xnor2_1 c665 (.A(net922),
    .B(net1078),
    .Y(net626));
 sky130_fd_sc_hd__clkbuf_2 c666 (.A(net728),
    .X(net627));
 sky130_fd_sc_hd__buf_1 c667 (.A(net728),
    .X(net628));
 sky130_fd_sc_hd__xnor2_1 c668 (.A(net517),
    .B(net625),
    .Y(net629));
 sky130_fd_sc_hd__xnor2_4 c669 (.A(net627),
    .B(net511),
    .Y(net630));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net988),
    .B(net27),
    .Y(net42));
 sky130_fd_sc_hd__a21bo_1 c670 (.A1(net630),
    .A2(net625),
    .B1_N(net996),
    .X(net631));
 sky130_fd_sc_hd__xnor2_1 c671 (.A(net621),
    .B(net630),
    .Y(net632));
 sky130_fd_sc_hd__a21bo_1 c672 (.A1(net508),
    .A2(net996),
    .B1_N(net625),
    .X(net633));
 sky130_fd_sc_hd__a21bo_2 c673 (.A1(net512),
    .A2(net109),
    .B1_N(net630),
    .X(net634));
 sky130_fd_sc_hd__xnor2_2 c674 (.A(net624),
    .B(net625),
    .Y(net635));
 sky130_fd_sc_hd__a31o_1 c675 (.A1(net632),
    .A2(net635),
    .A3(net996),
    .B1(net625),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net625),
    .A1(net634),
    .A2(net971),
    .A3(net622),
    .S0(net630),
    .S1(net996),
    .X(net637));
 sky130_fd_sc_hd__a41o_1 c677 (.A1(net526),
    .A2(net518),
    .A3(net634),
    .A4(net996),
    .B1(net630),
    .X(net638));
 sky130_fd_sc_hd__a41o_1 c678 (.A1(net511),
    .A2(net638),
    .A3(net528),
    .A4(net630),
    .B1(net996),
    .X(net639));
 sky130_fd_sc_hd__a31o_2 c679 (.A1(net635),
    .A2(net634),
    .A3(net971),
    .B1(net883),
    .X(net640));
 sky130_fd_sc_hd__a21bo_4 c68 (.A1(net1036),
    .A2(net41),
    .B1_N(net1016),
    .X(net43));
 sky130_fd_sc_hd__a41o_1 c680 (.A1(net630),
    .A2(net640),
    .A3(net250),
    .A4(net996),
    .B1(net1068),
    .X(net641));
 sky130_fd_sc_hd__xnor2_1 c681 (.A(net633),
    .B(net634),
    .Y(net642));
 sky130_fd_sc_hd__a41o_1 c682 (.A1(net138),
    .A2(net10),
    .A3(net635),
    .A4(net531),
    .B1(net875),
    .X(net643));
 sky130_fd_sc_hd__a21bo_1 c683 (.A1(net394),
    .A2(net539),
    .B1_N(net635),
    .X(net644));
 sky130_fd_sc_hd__a41o_1 c684 (.A1(net518),
    .A2(net528),
    .A3(net631),
    .A4(net873),
    .B1(net1064),
    .X(net645));
 sky130_fd_sc_hd__a21bo_1 c685 (.A1(net541),
    .A2(net987),
    .B1_N(net812),
    .X(net646));
 sky130_fd_sc_hd__a21bo_1 c686 (.A1(net398),
    .A2(net518),
    .B1_N(net376),
    .X(net647));
 sky130_fd_sc_hd__buf_1 c687 (.A(net918),
    .X(net648));
 sky130_fd_sc_hd__buf_1 c688 (.A(net915),
    .X(net649));
 sky130_fd_sc_hd__a21bo_1 c689 (.A1(net548),
    .A2(net634),
    .B1_N(net794),
    .X(net650));
 sky130_fd_sc_hd__xnor2_4 c69 (.A(net19),
    .B(net43),
    .Y(net44));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net635),
    .A1(net528),
    .A2(net539),
    .A3(net638),
    .S0(net647),
    .S1(net531),
    .X(net651));
 sky130_fd_sc_hd__buf_1 c691 (.A(net731),
    .X(net652));
 sky130_fd_sc_hd__a21bo_1 c692 (.A1(net629),
    .A2(net400),
    .B1_N(net649),
    .X(net653));
 sky130_fd_sc_hd__a21bo_1 c693 (.A1(net402),
    .A2(net539),
    .B1_N(net646),
    .X(net654));
 sky130_fd_sc_hd__dlymetal6s2s_1 c694 (.A(net920),
    .X(net655));
 sky130_fd_sc_hd__a21bo_1 c695 (.A1(net631),
    .A2(net652),
    .B1_N(net541),
    .X(net656));
 sky130_fd_sc_hd__a21bo_1 c696 (.A1(net376),
    .A2(net394),
    .B1_N(net959),
    .X(net657));
 sky130_fd_sc_hd__xnor2_2 c697 (.A(net648),
    .B(net656),
    .Y(net658));
 sky130_fd_sc_hd__a21bo_1 c698 (.A1(net657),
    .A2(net1060),
    .B1_N(net541),
    .X(net659));
 sky130_fd_sc_hd__a41o_2 c699 (.A1(net638),
    .A2(net394),
    .A3(net541),
    .A4(net623),
    .B1(net794),
    .X(net660));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net28),
    .B(net32),
    .Y(net45));
 sky130_fd_sc_hd__clkbuf_1 c700 (.A(net731),
    .X(net661));
 sky130_fd_sc_hd__xnor2_4 c701 (.A(net658),
    .B(net650),
    .Y(net662));
 sky130_fd_sc_hd__buf_1 c702 (.A(net806),
    .X(net663));
 sky130_fd_sc_hd__a21bo_1 c703 (.A1(net652),
    .A2(net661),
    .B1_N(net531),
    .X(net664));
 sky130_fd_sc_hd__a31o_1 c704 (.A1(net655),
    .A2(net518),
    .A3(net646),
    .B1(net559),
    .X(net665));
 sky130_fd_sc_hd__a31o_1 c705 (.A1(net665),
    .A2(net985),
    .A3(net569),
    .B1(net811),
    .X(net666));
 sky130_fd_sc_hd__a31o_1 c706 (.A1(net664),
    .A2(net418),
    .A3(net996),
    .B1(net634),
    .X(net667));
 sky130_fd_sc_hd__a31o_1 c707 (.A1(net655),
    .A2(net564),
    .A3(net569),
    .X(net809));
 sky130_fd_sc_hd__sdfbbp_1 c708 (.CLK(clknet_4_0_0_clk),
    .D(net666),
    .RESET_B(net660),
    .SCD(net998),
    .SCE(net664),
    .SET_B(net809),
    .Q(net670),
    .Q_N(net669));
 sky130_fd_sc_hd__sdfbbn_1 c709 (.CLK_N(clknet_4_0_0_clk),
    .D(net564),
    .RESET_B(net643),
    .SCD(net985),
    .SCE(net655),
    .SET_B(net1004),
    .Q(net671));
 sky130_fd_sc_hd__a21bo_4 c71 (.A1(net923),
    .A2(net27),
    .B1_N(net988),
    .X(net46));
 sky130_fd_sc_hd__buf_1 c710 (.A(net746),
    .X(net672));
 sky130_fd_sc_hd__sedfxbp_1 c711 (.CLK(clknet_4_0_0_clk),
    .D(net531),
    .DE(net564),
    .SCD(net664),
    .SCE(net660),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__sedfxbp_1 c712 (.CLK(clknet_4_0_0_clk),
    .D(net640),
    .DE(net671),
    .SCD(net548),
    .SCE(net660),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__buf_1 c713 (.A(net745),
    .X(net677));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net661),
    .A1(net663),
    .A2(net569),
    .A3(net998),
    .S0(net987),
    .S1(net873),
    .X(net678));
 sky130_fd_sc_hd__a21bo_1 c715 (.A1(net646),
    .A2(net30),
    .B1_N(clknet_1_0__leaf_net884),
    .X(net679));
 sky130_fd_sc_hd__a21bo_1 c716 (.A1(net649),
    .A2(net663),
    .B1_N(clknet_1_0__leaf_net884),
    .X(net680));
 sky130_fd_sc_hd__a31o_1 c717 (.A1(net674),
    .A2(net531),
    .A3(net646),
    .B1(clknet_1_0__leaf_net679),
    .X(net681));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(clknet_1_0__leaf_net680),
    .A1(net664),
    .A2(clknet_1_0__leaf_net679),
    .A3(net570),
    .S0(net873),
    .S1(net875),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net660),
    .A1(net649),
    .A2(net564),
    .A3(clknet_1_0__leaf_net679),
    .S0(net996),
    .S1(net640),
    .X(net683));
 sky130_fd_sc_hd__xnor2_1 c72 (.A(net40),
    .B(net44),
    .Y(net47));
 sky130_fd_sc_hd__buf_1 c720 (.A(net914),
    .X(net684));
 sky130_fd_sc_hd__sdfbbn_1 c721 (.CLK_N(clknet_4_0_0_clk),
    .D(net250),
    .RESET_B(net673),
    .SCD(net643),
    .SCE(clknet_1_0__leaf_net679),
    .SET_B(net660),
    .Q(net685));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net643),
    .A1(net649),
    .A2(net653),
    .A3(clknet_1_1__leaf_net680),
    .S0(net662),
    .S1(net787),
    .X(net686));
 sky130_fd_sc_hd__a31o_1 c723 (.A1(net685),
    .A2(net663),
    .A3(net998),
    .B1(clknet_1_0__leaf_net679),
    .X(net687));
 sky130_fd_sc_hd__a31o_1 c724 (.A1(net623),
    .A2(net687),
    .A3(net676),
    .B1(clknet_1_0__leaf_net679),
    .X(net688));
 sky130_fd_sc_hd__sedfxtp_1 c725 (.CLK(clknet_4_2_0_clk),
    .D(net688),
    .DE(net684),
    .SCD(clknet_1_1__leaf_net679),
    .SCE(net887),
    .Q(net689));
 sky130_fd_sc_hd__a41o_1 c726 (.A1(net123),
    .A2(clknet_1_1__leaf_net681),
    .A3(net999),
    .A4(net593),
    .B1(clknet_1_1__leaf_net884),
    .X(net690));
 sky130_fd_sc_hd__a41o_2 c727 (.A1(net937),
    .A2(net559),
    .A3(net123),
    .A4(net999),
    .B1(net787),
    .X(net691));
 sky130_fd_sc_hd__a31o_1 c728 (.A1(net556),
    .A2(net672),
    .A3(net548),
    .B1(clknet_1_0__leaf_net314),
    .X(net692));
 sky130_fd_sc_hd__sdfbbp_1 c729 (.CLK(clknet_4_2_0_clk),
    .D(net672),
    .RESET_B(clknet_1_0__leaf_net462),
    .SCD(net999),
    .SCE(net990),
    .SET_B(net874),
    .Q(net693));
 sky130_fd_sc_hd__a41o_2 c73 (.A1(net936),
    .A2(net45),
    .A3(net19),
    .A4(net42),
    .B1(net43),
    .X(net48));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net636),
    .A1(clknet_1_0__leaf_net595),
    .A2(net23),
    .A3(net593),
    .S0(net662),
    .S1(net691),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net684),
    .A1(clknet_1_1__leaf_net582),
    .A2(net515),
    .A3(net662),
    .S0(net787),
    .S1(net845),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net539),
    .A1(net694),
    .A2(net998),
    .A3(net626),
    .S0(clknet_1_0__leaf_net695),
    .S1(clknet_1_1__leaf_net885),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net670),
    .A1(net999),
    .A2(net678),
    .A3(net691),
    .S0(net593),
    .S1(clknet_1_1__leaf_net884),
    .X(net697));
 sky130_fd_sc_hd__sdfbbn_1 c734 (.CLK_N(clknet_4_2_0_clk),
    .D(net593),
    .RESET_B(net111),
    .SCD(net528),
    .SCE(net984),
    .SET_B(net691),
    .Q(net698));
 sky130_fd_sc_hd__a41o_1 c735 (.A1(net653),
    .A2(clknet_1_1__leaf_net695),
    .A3(clknet_1_1__leaf_net679),
    .A4(net266),
    .B1(net889),
    .X(net699));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net559),
    .A1(net697),
    .A2(net959),
    .A3(net677),
    .S0(net691),
    .S1(net937),
    .X(net700));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(clknet_1_0__leaf_net582),
    .A1(net548),
    .A2(net669),
    .A3(net691),
    .S0(net636),
    .S1(net889),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_0__leaf_net681),
    .A1(net266),
    .A2(net999),
    .A3(net971),
    .S0(net962),
    .S1(net874),
    .X(net702));
 sky130_fd_sc_hd__a41o_1 c739 (.A1(net701),
    .A2(net691),
    .A3(net983),
    .A4(net1004),
    .B1(clknet_1_1__leaf_net886),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 c74 (.A(net795),
    .X(net49));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net528),
    .A1(net698),
    .A2(net576),
    .A3(net266),
    .S0(net579),
    .S1(net889),
    .X(net704));
 sky130_fd_sc_hd__a31o_1 c741 (.A1(net983),
    .A2(net593),
    .A3(net691),
    .B1(clknet_1_0__leaf_net886),
    .X(net705));
 sky130_fd_sc_hd__a41o_1 c742 (.A1(net998),
    .A2(net691),
    .A3(net662),
    .A4(clknet_1_1__leaf_net679),
    .B1(net889),
    .X(net706));
 sky130_fd_sc_hd__sdfbbn_1 c743 (.CLK_N(clknet_4_2_0_clk),
    .D(net678),
    .RESET_B(net703),
    .SCD(net705),
    .SCE(net691),
    .SET_B(net515),
    .Q(net707));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net634),
    .A1(clknet_1_0__leaf_net695),
    .A2(net548),
    .A3(net691),
    .S0(net844),
    .S1(clknet_1_0__leaf_net885),
    .X(net708));
 sky130_fd_sc_hd__a41o_1 c745 (.A1(net700),
    .A2(clknet_1_1__leaf_net595),
    .A3(net111),
    .A4(net891),
    .B1(net893),
    .X(net709));
 sky130_fd_sc_hd__sdfbbp_1 c746 (.CLK(clknet_4_2_0_clk),
    .D(net626),
    .RESET_B(net944),
    .SCD(net30),
    .SCE(net797),
    .SET_B(net892),
    .Q(net710));
 sky130_fd_sc_hd__a41o_1 c747 (.A1(net707),
    .A2(net709),
    .A3(net710),
    .A4(net573),
    .B1(net890),
    .X(net711));
 sky130_fd_sc_hd__mux4_2 c748 (.A0(net215),
    .A1(net612),
    .A2(net30),
    .A3(net888),
    .S0(net890),
    .S1(net893),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net579),
    .A1(net612),
    .A2(net712),
    .A3(net925),
    .S0(net215),
    .S1(clknet_1_0__leaf_net473),
    .X(net713));
 sky130_fd_sc_hd__xnor2_2 c75 (.A(net8),
    .B(net49),
    .Y(net50));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net266),
    .A1(net569),
    .A2(net689),
    .A3(net1023),
    .S0(net867),
    .S1(net890),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net677),
    .A1(net1023),
    .A2(clknet_1_0__leaf_net473),
    .A3(clknet_1_1__leaf_net679),
    .S0(net1004),
    .S1(net893),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net602),
    .A1(net1015),
    .A2(net607),
    .A3(net867),
    .S0(net882),
    .S1(net893),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_1__leaf_net679),
    .A1(net471),
    .A2(net215),
    .A3(net609),
    .S0(net569),
    .S1(net882),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net706),
    .A1(net570),
    .A2(net30),
    .A3(net712),
    .S0(net867),
    .S1(net882),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net628),
    .A1(net715),
    .A2(net714),
    .A3(clknet_1_0__leaf_net473),
    .S0(net570),
    .S1(net893),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net662),
    .A1(net1013),
    .A2(clknet_1_1__leaf_net679),
    .A3(net1025),
    .S0(net815),
    .S1(net890),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net689),
    .A1(net576),
    .A2(clknet_1_0__leaf_net473),
    .A3(net1004),
    .S0(net882),
    .S1(net894),
    .X(net721));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net608),
    .A1(net569),
    .A2(net718),
    .A3(net570),
    .S0(net662),
    .S1(net893),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net1015),
    .A1(clknet_1_0__leaf_net314),
    .A2(net711),
    .A3(net609),
    .S0(net1024),
    .S1(net895),
    .X(net723));
 sky130_fd_sc_hd__a21bo_4 c76 (.A1(net930),
    .A2(net50),
    .B1_N(net1033),
    .X(net51));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net693),
    .A1(clknet_1_1__leaf_net462),
    .A2(net717),
    .A3(net30),
    .S0(net895),
    .S1(net896),
    .X(net724));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net721),
    .A1(net798),
    .A2(net882),
    .A3(net893),
    .S0(net895),
    .S1(net897),
    .X(net725));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net609),
    .A1(net716),
    .A2(net720),
    .A3(net725),
    .S0(net1026),
    .S1(net896),
    .X(net726));
 sky130_fd_sc_hd__xnor2_1 c77 (.A(net931),
    .B(net31),
    .Y(net52));
 sky130_fd_sc_hd__a21bo_4 c78 (.A1(net11),
    .A2(net988),
    .B1_N(net926),
    .X(net967));
 sky130_fd_sc_hd__a31o_2 c79 (.A1(net989),
    .A2(net49),
    .A3(net52),
    .B1(net41),
    .X(net53));
 sky130_fd_sc_hd__xnor2_4 c80 (.A(net1017),
    .B(net992),
    .Y(net948));
 sky130_fd_sc_hd__xnor2_4 c81 (.A(net53),
    .B(net43),
    .Y(net54));
 sky130_fd_sc_hd__xnor2_2 c82 (.A(net13),
    .B(net988),
    .Y(net55));
 sky130_fd_sc_hd__a41o_1 c83 (.A1(net37),
    .A2(net48),
    .A3(net45),
    .A4(net1034),
    .B1(net44),
    .X(net56));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net44),
    .A1(net48),
    .A2(net51),
    .A3(net50),
    .S0(net989),
    .S1(net55),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net46),
    .A1(net56),
    .A2(net55),
    .A3(net57),
    .S0(net989),
    .S1(net1035),
    .X(net58));
 sky130_fd_sc_hd__buf_1 c86 (.A(net795),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net43),
    .A1(net53),
    .A2(net59),
    .A3(net57),
    .S0(net1037),
    .S1(net51),
    .X(net60));
 sky130_fd_sc_hd__xnor2_1 c88 (.A(net3),
    .B(net13),
    .Y(net61));
 sky130_fd_sc_hd__xnor2_1 c89 (.A(net3),
    .B(net54),
    .Y(net62));
 sky130_fd_sc_hd__xnor2_1 c90 (.A(net52),
    .B(net42),
    .Y(net63));
 sky130_fd_sc_hd__a21bo_1 c91 (.A1(net61),
    .A2(net41),
    .B1_N(net973),
    .X(net64));
 sky130_fd_sc_hd__xnor2_1 c92 (.A(net940),
    .B(net23),
    .Y(net65));
 sky130_fd_sc_hd__xnor2_1 c93 (.A(net64),
    .B(net24),
    .Y(net66));
 sky130_fd_sc_hd__mux4_1 c94 (.A0(net66),
    .A1(net3),
    .A2(net13),
    .A3(net45),
    .S0(net19),
    .S1(net948),
    .X(net67));
 sky130_fd_sc_hd__xnor2_1 c95 (.A(net41),
    .B(net51),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_1 c96 (.A(net53),
    .B(net973),
    .Y(net69));
 sky130_fd_sc_hd__buf_1 c97 (.A(net810),
    .X(net70));
 sky130_fd_sc_hd__a21bo_1 c98 (.A1(net944),
    .A2(net48),
    .B1_N(net972),
    .X(net71));
 sky130_fd_sc_hd__xnor2_1 c99 (.A(net68),
    .B(net13),
    .Y(net72));
 sky130_fd_sc_hd__mux4_1 merge763 (.A0(net47),
    .A1(net43),
    .A2(net57),
    .A3(net52),
    .S0(net45),
    .S1(net822),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_1 merge764 (.A(net919),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 merge765 (.A(net915),
    .X(net729));
 sky130_fd_sc_hd__buf_1 merge766 (.A(clknet_1_1__leaf_net905),
    .X(net730));
 sky130_fd_sc_hd__sedfxtp_1 merge767 (.CLK(clknet_4_1_0_clk),
    .D(net642),
    .DE(net398),
    .SCD(net400),
    .SCE(net657),
    .Q(net731));
 sky130_fd_sc_hd__sedfxtp_1 merge768 (.CLK(clknet_4_13_0_clk),
    .D(net89),
    .DE(net84),
    .SCD(net92),
    .SCE(net1069),
    .Q(net732));
 sky130_fd_sc_hd__a31o_1 merge769 (.A1(net1038),
    .A2(net56),
    .A3(net47),
    .B1(net26),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net970),
    .A1(clknet_1_0__leaf_net456),
    .A2(net111),
    .A3(clknet_1_0__leaf_net464),
    .S0(net844),
    .S1(net861),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_1 merge771 (.A(net778),
    .X(net735));
 sky130_fd_sc_hd__a31o_1 merge772 (.A1(net941),
    .A2(net150),
    .A3(net133),
    .B1(net147),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net419),
    .A1(net984),
    .A2(net970),
    .A3(clknet_1_1__leaf_net411),
    .S0(net420),
    .S1(net422),
    .X(net737));
 sky130_fd_sc_hd__buf_1 merge774 (.A(clknet_1_0__leaf_net905),
    .X(net738));
 sky130_fd_sc_hd__a31o_1 merge775 (.A1(net399),
    .A2(net389),
    .A3(net378),
    .B1(clknet_1_0__leaf_net964),
    .X(net739));
 sky130_fd_sc_hd__sdfrbp_1 merge776 (.CLK(clknet_4_12_0_clk),
    .D(net190),
    .RESET_B(net57),
    .SCD(net268),
    .SCE(net152),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__a41o_1 merge777 (.A1(net82),
    .A2(net170),
    .A3(net191),
    .A4(net197),
    .B1(net173),
    .X(net742));
 sky130_fd_sc_hd__sdfrbp_1 merge778 (.CLK(clknet_4_1_0_clk),
    .D(net551),
    .RESET_B(net424),
    .SCD(net534),
    .SCE(net557),
    .Q(net744),
    .Q_N(net743));
 sky130_fd_sc_hd__sdfbbn_1 merge779 (.CLK_N(clknet_4_0_0_clk),
    .D(net417),
    .RESET_B(net640),
    .SCD(net998),
    .SCE(net675),
    .SET_B(net655),
    .Q(net746),
    .Q_N(net745));
 sky130_fd_sc_hd__a41o_1 merge780 (.A1(net143),
    .A2(net986),
    .A3(net141),
    .A4(net977),
    .B1(net131),
    .X(net747));
 sky130_fd_sc_hd__a41o_1 merge781 (.A1(net175),
    .A2(net50),
    .A3(net1006),
    .A4(net183),
    .B1(net8),
    .X(net748));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net553),
    .A1(net448),
    .A2(net550),
    .A3(net575),
    .S0(net574),
    .S1(clknet_1_0__leaf_net314),
    .X(net749));
 sky130_fd_sc_hd__sdfrtn_1 merge783 (.CLK_N(clknet_4_9_0_clk),
    .D(net1058),
    .RESET_B(net480),
    .SCD(net409),
    .SCE(net214),
    .Q(net750));
 sky130_fd_sc_hd__clkbuf_1 merge784 (.A(net917),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net481),
    .A1(net471),
    .A2(net336),
    .A3(net330),
    .S0(net78),
    .S1(net833),
    .X(net752));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net550),
    .A1(net555),
    .A2(net484),
    .A3(net476),
    .S0(net992),
    .S1(net844),
    .X(net753));
 sky130_fd_sc_hd__a41o_1 merge787 (.A1(net407),
    .A2(net1055),
    .A3(net378),
    .A4(net959),
    .B1(net927),
    .X(net754));
 sky130_fd_sc_hd__sdfbbn_1 merge788 (.CLK_N(clknet_4_13_0_clk),
    .D(net56),
    .RESET_B(net71),
    .SCD(net154),
    .SCE(net152),
    .SET_B(net968),
    .Q(net756),
    .Q_N(net755));
 sky130_fd_sc_hd__a31o_1 merge789 (.A1(net391),
    .A2(net510),
    .A3(net513),
    .B1(net516),
    .X(net757));
 sky130_fd_sc_hd__a31o_1 merge790 (.A1(net293),
    .A2(net292),
    .A3(net294),
    .B1(clknet_1_0__leaf_net290),
    .X(net758));
 sky130_fd_sc_hd__sdfbbp_1 merge791 (.CLK(clknet_4_9_0_clk),
    .D(net460),
    .RESET_B(net469),
    .SCD(net342),
    .SCE(net466),
    .SET_B(net214),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__sdfrtp_1 merge792 (.CLK(clknet_4_12_0_clk),
    .D(net307),
    .RESET_B(net292),
    .SCD(net321),
    .SCE(net317),
    .Q(net761));
 sky130_fd_sc_hd__sdfbbn_1 merge793 (.CLK_N(clknet_4_5_0_clk),
    .D(net288),
    .RESET_B(net155),
    .SCD(net256),
    .SCE(net141),
    .SET_B(net268),
    .Q(net763),
    .Q_N(net762));
 sky130_fd_sc_hd__sdfbbn_1 merge794 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net309),
    .RESET_B(net307),
    .SCD(net18),
    .SCE(net39),
    .SET_B(net152),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__a31o_1 merge795 (.A1(net521),
    .A2(net516),
    .A3(net1000),
    .B1(net536),
    .X(net766));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net583),
    .A1(net515),
    .A2(net389),
    .A3(net178),
    .S0(clknet_1_0__leaf_net462),
    .S1(net864),
    .X(net767));
 sky130_fd_sc_hd__mux4_1 merge797 (.A0(net532),
    .A1(net533),
    .A2(clknet_1_0__leaf_net964),
    .A3(net1062),
    .S0(net660),
    .S1(net656),
    .X(net768));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net155),
    .A1(net283),
    .A2(net286),
    .A3(net268),
    .S0(net239),
    .S1(net261),
    .X(net769));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net199),
    .A1(net82),
    .A2(net198),
    .A3(net160),
    .S0(net205),
    .S1(net191),
    .X(net770));
 sky130_fd_sc_hd__mux4_1 merge800 (.A0(net308),
    .A1(net319),
    .A2(net54),
    .A3(net92),
    .S0(net972),
    .S1(net807),
    .X(net771));
 sky130_fd_sc_hd__mux4_1 merge801 (.A0(net62),
    .A1(net73),
    .A2(net972),
    .A3(net97),
    .S0(net95),
    .S1(net96),
    .X(net772));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net516),
    .A1(net396),
    .A2(net518),
    .A3(net520),
    .S0(net940),
    .S1(net519),
    .X(net773));
 sky130_fd_sc_hd__mux4_1 merge803 (.A0(net39),
    .A1(net133),
    .A2(net571),
    .A3(net783),
    .S0(net787),
    .S1(net876),
    .X(net774));
 sky130_fd_sc_hd__mux4_1 merge804 (.A0(net545),
    .A1(net531),
    .A2(net536),
    .A3(net444),
    .S0(net996),
    .S1(clknet_1_0__leaf_net679),
    .X(net775));
 sky130_fd_sc_hd__mux4_1 merge805 (.A0(net644),
    .A1(net640),
    .A2(net932),
    .A3(net510),
    .S0(net976),
    .S1(net873),
    .X(net776));
 sky130_fd_sc_hd__mux4_1 merge806 (.A0(net554),
    .A1(net543),
    .A2(net557),
    .A3(net540),
    .S0(net537),
    .S1(net528),
    .X(net777));
 sky130_fd_sc_hd__sdfbbp_1 merge807 (.CLK(clknet_4_1_0_clk),
    .D(net537),
    .RESET_B(net543),
    .SCD(net536),
    .SCE(net509),
    .SET_B(net535),
    .Q(net779),
    .Q_N(net778));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net541),
    .A1(net644),
    .A2(net647),
    .A3(net110),
    .S0(net378),
    .S1(net259),
    .X(net780));
 sky130_fd_sc_hd__mux4_1 merge809 (.A0(net647),
    .A1(net654),
    .A2(net622),
    .A3(net257),
    .S0(net108),
    .S1(net874),
    .X(net781));
 sky130_fd_sc_hd__dfrbp_1 merge810 (.CLK(clknet_4_3_0_clk),
    .D(net588),
    .RESET_B(net592),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dfrbp_1 merge811 (.CLK(clknet_4_14_0_clk),
    .D(net352),
    .RESET_B(net356),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dfrtn_1 merge812 (.CLK_N(clknet_4_13_0_clk),
    .D(net211),
    .RESET_B(net742),
    .Q(net786));
 sky130_fd_sc_hd__dfrtp_1 merge813 (.CLK(clknet_4_5_0_clk),
    .D(net280),
    .Q(net281));
 sky130_fd_sc_hd__dfrtp_1 merge814 (.CLK(clknet_4_15_0_clk),
    .D(net86),
    .RESET_B(net105),
    .Q(net788));
 sky130_fd_sc_hd__dfrtp_1 merge815 (.CLK(clknet_4_11_0_clk),
    .D(net507),
    .RESET_B(net493),
    .Q(net789));
 sky130_fd_sc_hd__dfsbp_2 merge816 (.CLK(clknet_4_7_0_clk),
    .D(net167),
    .SET_B(net736),
    .Q(net791),
    .Q_N(net790));
 sky130_fd_sc_hd__dfsbp_1 merge817 (.CLK(clknet_4_3_0_clk),
    .D(net558),
    .SET_B(net567),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__dfstp_1 merge818 (.CLK(clknet_4_0_0_clk),
    .D(net645),
    .SET_B(net659),
    .Q(net794));
 sky130_fd_sc_hd__dfstp_2 merge819 (.CLK(clknet_4_13_0_clk),
    .D(net727),
    .SET_B(net60),
    .Q(net795));
 sky130_fd_sc_hd__dfstp_1 merge820 (.CLK(clknet_4_5_0_clk),
    .D(net739),
    .SET_B(net754),
    .Q(net796));
 sky130_fd_sc_hd__dlrbn_1 merge821 (.D(net690),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net692),
    .Q(net798),
    .Q_N(net797));
 sky130_fd_sc_hd__dlrbn_1 merge822 (.D(net757),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net766),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlrbp_1 merge823 (.D(net452),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net463),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dlrbp_1 merge824 (.D(net234),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net233),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlrtn_1 merge825 (.D(net334),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net337),
    .Q(net805));
 sky130_fd_sc_hd__dlrtn_1 merge826 (.D(net546),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net768),
    .Q(net806));
 sky130_fd_sc_hd__dlrtn_1 merge827 (.D(net325),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net316),
    .Q(net807));
 sky130_fd_sc_hd__dlrtp_1 merge828 (.D(net599),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net614),
    .Q(net808));
 sky130_fd_sc_hd__dlrtp_1 merge829 (.D(net667),
    .GATE(clknet_4_0_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dlrtp_1 merge830 (.D(net76),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net733),
    .Q(net810));
 sky130_fd_sc_hd__edfxbp_1 merge831 (.CLK(clknet_4_0_0_clk),
    .D(net639),
    .DE(net641),
    .Q(net812),
    .Q_N(net811));
 sky130_fd_sc_hd__edfxtp_1 merge832 (.CLK(clknet_4_7_0_clk),
    .D(net748),
    .DE(net172),
    .Q(net813));
 sky130_fd_sc_hd__sdlclkp_1 merge833 (.CLK(clknet_4_7_0_clk),
    .GATE(net297),
    .SCE(net758),
    .GCLK(net814));
 sky130_fd_sc_hd__sdlclkp_2 merge834 (.CLK(clknet_4_8_0_clk),
    .GATE(net726),
    .SCE(net713),
    .GCLK(net815));
 sky130_fd_sc_hd__sdlclkp_4 merge835 (.CLK(clknet_4_6_0_clk),
    .GATE(net434),
    .SCE(net435),
    .GCLK(net816));
 sky130_fd_sc_hd__dfrbp_2 merge836 (.CLK(clknet_4_5_0_clk),
    .D(net392),
    .RESET_B(net395),
    .Q(net818),
    .Q_N(net817));
 sky130_fd_sc_hd__dfrbp_1 merge837 (.CLK(clknet_4_8_0_clk),
    .D(net478),
    .RESET_B(net487),
    .Q(net820),
    .Q_N(net819));
 sky130_fd_sc_hd__dfrtn_1 merge838 (.CLK_N(clknet_4_10_0_clk),
    .D(net699),
    .RESET_B(net506),
    .Q(net962));
 sky130_fd_sc_hd__dfrtp_2 merge839 (.CLK(clknet_4_3_0_clk),
    .D(net438),
    .RESET_B(net572),
    .Q(net946));
 sky130_fd_sc_hd__dfrtp_4 merge840 (.CLK(clknet_4_5_0_clk),
    .D(net747),
    .RESET_B(net156),
    .Q(net821));
 sky130_fd_sc_hd__dfxbp_2 s841 (.CLK(clknet_4_13_0_clk),
    .D(net58),
    .Q(net823),
    .Q_N(net822));
 sky130_fd_sc_hd__dfxbp_1 s842 (.CLK(clknet_4_13_0_clk),
    .D(net67),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dfxtp_1 s843 (.CLK(clknet_4_13_0_clk),
    .D(net81),
    .Q(net826));
 sky130_fd_sc_hd__dfxtp_1 s844 (.CLK(clknet_4_13_0_clk),
    .D(net83),
    .Q(net827));
 sky130_fd_sc_hd__dfxtp_2 s845 (.CLK(clknet_4_15_0_clk),
    .D(net102),
    .Q(net950));
 sky130_fd_sc_hd__dlclkp_1 s846 (.CLK(clknet_4_15_0_clk),
    .GATE(net104),
    .GCLK(net828));
 sky130_fd_sc_hd__dlclkp_2 s847 (.CLK(clknet_4_15_0_clk),
    .GATE(net106),
    .GCLK(net829));
 sky130_fd_sc_hd__dlclkp_4 s848 (.CLK(clknet_4_15_0_clk),
    .GATE(net107),
    .GCLK(net830));
 sky130_fd_sc_hd__dlxbn_1 s849 (.D(net212),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net832),
    .Q_N(net831));
 sky130_fd_sc_hd__dlxbn_1 s850 (.D(net213),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net834),
    .Q_N(net833));
 sky130_fd_sc_hd__dlxbp_1 s851 (.D(net228),
    .GATE(clknet_4_15_0_clk),
    .Q(net836),
    .Q_N(net835));
 sky130_fd_sc_hd__dlxtn_1 s852 (.D(net235),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net837));
 sky130_fd_sc_hd__dlxtn_1 s853 (.D(net236),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net838));
 sky130_fd_sc_hd__dlxtn_2 s854 (.D(net299),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net839));
 sky130_fd_sc_hd__dlxtp_1 s855 (.D(net301),
    .GATE(clknet_4_7_0_clk),
    .Q(net840));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s856 (.D(net302),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net841));
 sky130_fd_sc_hd__dfxbp_1 s857 (.CLK(clknet_4_12_0_clk),
    .D(net323),
    .Q(net843),
    .Q_N(net842));
 sky130_fd_sc_hd__dfxbp_1 s858 (.CLK(clknet_4_9_0_clk),
    .D(net324),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__dfxtp_1 s859 (.CLK(clknet_4_9_0_clk),
    .D(net344),
    .Q(net846));
 sky130_fd_sc_hd__dfxtp_1 s860 (.CLK(clknet_4_14_0_clk),
    .D(net349),
    .Q(net847));
 sky130_fd_sc_hd__dfxtp_1 s861 (.CLK(clknet_4_15_0_clk),
    .D(net360),
    .Q(net848));
 sky130_fd_sc_hd__dlclkp_1 s862 (.CLK(clknet_4_14_0_clk),
    .GATE(net367),
    .GCLK(net849));
 sky130_fd_sc_hd__dlclkp_2 s863 (.CLK(clknet_4_14_0_clk),
    .GATE(net370),
    .GCLK(net850));
 sky130_fd_sc_hd__dlclkp_4 s864 (.CLK(clknet_4_14_0_clk),
    .GATE(net371),
    .GCLK(net851));
 sky130_fd_sc_hd__dlxbn_1 s865 (.D(net374),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net853),
    .Q_N(net852));
 sky130_fd_sc_hd__dlxbn_1 s866 (.D(net416),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net855),
    .Q_N(net854));
 sky130_fd_sc_hd__dlxbp_1 s867 (.D(net429),
    .GATE(clknet_4_4_0_clk),
    .Q(net857),
    .Q_N(net856));
 sky130_fd_sc_hd__dlxtn_1 s868 (.D(net437),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net858));
 sky130_fd_sc_hd__dlxtn_1 s869 (.D(net440),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net859));
 sky130_fd_sc_hd__dlxtn_1 s870 (.D(net442),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net860));
 sky130_fd_sc_hd__dlxtp_1 s871 (.D(net453),
    .GATE(clknet_4_6_0_clk),
    .Q(net861));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s872 (.D(net454),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net862));
 sky130_fd_sc_hd__dfxbp_1 s873 (.CLK(clknet_4_10_0_clk),
    .D(net465),
    .Q(net952),
    .Q_N(net863));
 sky130_fd_sc_hd__dfxbp_1 s874 (.CLK(clknet_4_3_0_clk),
    .D(net468),
    .Q(net865),
    .Q_N(net864));
 sky130_fd_sc_hd__dfxtp_1 s875 (.CLK(clknet_4_11_0_clk),
    .D(net470),
    .Q(net866));
 sky130_fd_sc_hd__dfxtp_2 s876 (.CLK(clknet_4_10_0_clk),
    .D(net485),
    .Q(net867));
 sky130_fd_sc_hd__dfxtp_1 s877 (.CLK(clknet_4_11_0_clk),
    .D(net490),
    .Q(net955));
 sky130_fd_sc_hd__dlclkp_1 s878 (.CLK(clknet_4_11_0_clk),
    .GATE(net494),
    .GCLK(net868));
 sky130_fd_sc_hd__dlclkp_2 s879 (.CLK(clknet_4_11_0_clk),
    .GATE(net495),
    .GCLK(net869));
 sky130_fd_sc_hd__dlclkp_4 s880 (.CLK(clknet_4_14_0_clk),
    .GATE(net496),
    .GCLK(net963));
 sky130_fd_sc_hd__dlxbn_1 s881 (.D(net500),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net870));
 sky130_fd_sc_hd__dlxbn_1 s882 (.D(net501),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net871));
 sky130_fd_sc_hd__dlxbp_1 s883 (.D(net503),
    .GATE(clknet_4_11_0_clk),
    .Q(net872));
 sky130_fd_sc_hd__dlxtn_1 s884 (.D(net504),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net961));
 sky130_fd_sc_hd__dlxtn_2 s885 (.D(net529),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net873));
 sky130_fd_sc_hd__dlxtn_2 s886 (.D(net544),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net874));
 sky130_fd_sc_hd__dlxtp_1 s887 (.D(net547),
    .GATE(clknet_4_1_0_clk),
    .Q(net875));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s888 (.D(net589),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dfxbp_1 s889 (.CLK(clknet_4_3_0_clk),
    .D(net594),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dfxbp_1 s890 (.CLK(clknet_4_8_0_clk),
    .D(net604),
    .Q(net880),
    .Q_N(net879));
 sky130_fd_sc_hd__dfxtp_1 s891 (.CLK(clknet_4_10_0_clk),
    .D(net618),
    .Q(net881));
 sky130_fd_sc_hd__dfxtp_2 s892 (.CLK(clknet_4_10_0_clk),
    .D(net620),
    .Q(net882));
 sky130_fd_sc_hd__dfxtp_1 s893 (.CLK(clknet_4_0_0_clk),
    .D(net637),
    .Q(net883));
 sky130_fd_sc_hd__dlclkp_1 s894 (.CLK(clknet_4_0_0_clk),
    .GATE(net651),
    .GCLK(net884));
 sky130_fd_sc_hd__dlclkp_2 s895 (.CLK(clknet_4_2_0_clk),
    .GATE(net682),
    .GCLK(net885));
 sky130_fd_sc_hd__dlclkp_4 s896 (.CLK(clknet_4_2_0_clk),
    .GATE(net683),
    .GCLK(net886));
 sky130_fd_sc_hd__dlxbn_1 s897 (.D(net686),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__dlxbn_1 s898 (.D(net696),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net890),
    .Q_N(net889));
 sky130_fd_sc_hd__dlxbp_1 s899 (.D(net702),
    .GATE(clknet_4_2_0_clk),
    .Q(net891));
 sky130_fd_sc_hd__dlxtn_1 s900 (.D(net704),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net892));
 sky130_fd_sc_hd__dlxtn_2 s901 (.D(net708),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net893));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net719),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net894));
 sky130_fd_sc_hd__dlxtp_1 s903 (.D(net722),
    .GATE(clknet_4_8_0_clk),
    .Q(net895));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s904 (.D(net723),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net896));
 sky130_fd_sc_hd__dfxbp_1 s905 (.CLK(clknet_4_10_0_clk),
    .D(net724),
    .Q(net897));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_4_6_0_clk),
    .D(net734),
    .Q(net899),
    .Q_N(net898));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_6_0_clk),
    .D(net737),
    .Q(net900));
 sky130_fd_sc_hd__dfxtp_1 s908 (.CLK(clknet_4_3_0_clk),
    .D(net749),
    .Q(net901));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_4_11_0_clk),
    .D(net752),
    .Q(net902));
 sky130_fd_sc_hd__dlclkp_1 s910 (.CLK(clknet_4_3_0_clk),
    .GATE(net753),
    .GCLK(net903));
 sky130_fd_sc_hd__dlclkp_2 s911 (.CLK(clknet_4_3_0_clk),
    .GATE(net767),
    .GCLK(net904));
 sky130_fd_sc_hd__dlclkp_4 s912 (.CLK(clknet_4_5_0_clk),
    .GATE(net769),
    .GCLK(net905));
 sky130_fd_sc_hd__dlxbn_1 s913 (.D(net770),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net907),
    .Q_N(net906));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net771),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net909),
    .Q_N(net908));
 sky130_fd_sc_hd__dlxbp_1 s915 (.D(net772),
    .GATE(clknet_4_13_0_clk),
    .Q(net911),
    .Q_N(net910));
 sky130_fd_sc_hd__dlxtn_1 s916 (.D(net773),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net912));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net774),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net913));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net775),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net914));
 sky130_fd_sc_hd__dlxtp_1 s919 (.D(net776),
    .GATE(clknet_4_1_0_clk),
    .Q(net915));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s920 (.D(net777),
    .SLEEP_B(clknet_4_1_0_clk),
    .Q(net916));
 sky130_fd_sc_hd__dfxbp_1 s921 (.CLK(clknet_4_4_0_clk),
    .D(net780),
    .Q(net918),
    .Q_N(net917));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_4_0_0_clk),
    .D(net781),
    .Q(net920),
    .Q_N(net919));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_8 input1 (.A(in0),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net922));
 sky130_fd_sc_hd__buf_6 input4 (.A(in11),
    .X(net923));
 sky130_fd_sc_hd__buf_2 input5 (.A(in12),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net925));
 sky130_fd_sc_hd__buf_4 input7 (.A(in14),
    .X(net926));
 sky130_fd_sc_hd__buf_4 input8 (.A(in15),
    .X(net927));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(in17),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net930));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(in19),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(in2),
    .X(net932));
 sky130_fd_sc_hd__buf_2 input14 (.A(in20),
    .X(net933));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net934));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net935));
 sky130_fd_sc_hd__buf_4 input17 (.A(in23),
    .X(net936));
 sky130_fd_sc_hd__buf_8 input18 (.A(in24),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in3),
    .X(net938));
 sky130_fd_sc_hd__buf_4 input20 (.A(in4),
    .X(net939));
 sky130_fd_sc_hd__buf_4 input21 (.A(in5),
    .X(net940));
 sky130_fd_sc_hd__buf_2 input22 (.A(in6),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(in7),
    .X(net942));
 sky130_fd_sc_hd__buf_4 input24 (.A(in8),
    .X(net943));
 sky130_fd_sc_hd__buf_2 input25 (.A(in9),
    .X(net944));
 sky130_fd_sc_hd__buf_2 output26 (.A(net945),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output27 (.A(net946),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net1031),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output29 (.A(net948),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output30 (.A(net949),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net950),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output32 (.A(net951),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output33 (.A(net952),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output34 (.A(net953),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output35 (.A(net954),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output36 (.A(net955),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output37 (.A(net956),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output38 (.A(net985),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net958),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output40 (.A(net959),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output41 (.A(net960),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output42 (.A(net961),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output43 (.A(net962),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(clknet_1_1__leaf_net963),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(clknet_1_0__leaf_net964),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output46 (.A(net987),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net966),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net967),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net980),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output50 (.A(net969),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net445),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_8 fanout52 (.A(net260),
    .X(net971));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net975),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(net975),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(net63),
    .X(net975));
 sky130_fd_sc_hd__buf_4 max_cap57 (.A(net380),
    .X(net976));
 sky130_fd_sc_hd__buf_4 max_cap58 (.A(net137),
    .X(net977));
 sky130_fd_sc_hd__buf_4 max_cap59 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__buf_4 max_cap60 (.A(net250),
    .X(net979));
 sky130_fd_sc_hd__buf_4 max_cap61 (.A(net968),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net84),
    .X(net981));
 sky130_fd_sc_hd__buf_6 wire63 (.A(net25),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net397),
    .X(net983));
 sky130_fd_sc_hd__buf_8 fanout65 (.A(net249),
    .X(net984));
 sky130_fd_sc_hd__buf_4 max_cap66 (.A(net957),
    .X(net985));
 sky130_fd_sc_hd__buf_4 max_cap67 (.A(net128),
    .X(net986));
 sky130_fd_sc_hd__buf_4 max_cap68 (.A(net965),
    .X(net987));
 sky130_fd_sc_hd__buf_4 max_cap69 (.A(net41),
    .X(net988));
 sky130_fd_sc_hd__buf_12 fanout70 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__buf_12 fanout71 (.A(net17),
    .X(net990));
 sky130_fd_sc_hd__buf_4 max_cap72 (.A(net125),
    .X(net991));
 sky130_fd_sc_hd__buf_4 max_cap73 (.A(net29),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net335),
    .X(net993));
 sky130_fd_sc_hd__buf_4 max_cap75 (.A(net269),
    .X(net994));
 sky130_fd_sc_hd__buf_4 max_cap76 (.A(net1022),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net628),
    .X(net996));
 sky130_fd_sc_hd__buf_4 max_cap78 (.A(net40),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(net439),
    .X(net998));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(net573),
    .X(net999));
 sky130_fd_sc_hd__buf_4 wire81 (.A(net246),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 max_cap82 (.A(net243),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net157),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 max_cap84 (.A(net114),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_8 fanout85 (.A(net839),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net221),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 max_cap87 (.A(net134),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 max_cap88 (.A(net115),
    .X(net1007));
 sky130_fd_sc_hd__buf_8 max_cap89 (.A(net111),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net905 (.A(net905),
    .X(clknet_0_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_0__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net905 (.A(clknet_0_net905),
    .X(clknet_1_1__leaf_net905));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net738 (.A(net738),
    .X(clknet_0_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_0__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net738 (.A(clknet_0_net738),
    .X(clknet_1_1__leaf_net738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net276 (.A(net276),
    .X(clknet_0_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_0__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net276 (.A(clknet_0_net276),
    .X(clknet_1_1__leaf_net276));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net279 (.A(net279),
    .X(clknet_0_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_0__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net279 (.A(clknet_0_net279),
    .X(clknet_1_1__leaf_net279));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net408 (.A(net408),
    .X(clknet_0_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_0__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net502 (.A(net502),
    .X(clknet_0_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_0__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net502 (.A(clknet_0_net502),
    .X(clknet_1_1__leaf_net502));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net964 (.A(net964),
    .X(clknet_0_net964));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net964 (.A(clknet_0_net964),
    .X(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net964 (.A(clknet_0_net964),
    .X(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net412 (.A(net412),
    .X(clknet_0_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_0__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net412 (.A(clknet_0_net412),
    .X(clknet_1_1__leaf_net412));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net410 (.A(net410),
    .X(clknet_0_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_0__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net410 (.A(clknet_0_net410),
    .X(clknet_1_1__leaf_net410));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net270 (.A(net270),
    .X(clknet_0_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_0__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net270 (.A(clknet_0_net270),
    .X(clknet_1_1__leaf_net270));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net273 (.A(net273),
    .X(clknet_0_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_0__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net273 (.A(clknet_0_net273),
    .X(clknet_1_1__leaf_net273));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net730 (.A(net730),
    .X(clknet_0_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net730 (.A(clknet_0_net730),
    .X(clknet_1_0__leaf_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net730 (.A(clknet_0_net730),
    .X(clknet_1_1__leaf_net730));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net814 (.A(net814),
    .X(clknet_0_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_0__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net814 (.A(clknet_0_net814),
    .X(clknet_1_1__leaf_net814));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net304 (.A(net304),
    .X(clknet_0_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net304 (.A(clknet_0_net304),
    .X(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net304 (.A(clknet_0_net304),
    .X(clknet_1_1__leaf_net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net473 (.A(net473),
    .X(clknet_0_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_0__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net473 (.A(clknet_0_net473),
    .X(clknet_1_1__leaf_net473));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net459 (.A(net459),
    .X(clknet_0_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_0__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net459 (.A(clknet_0_net459),
    .X(clknet_1_1__leaf_net459));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net464 (.A(net464),
    .X(clknet_0_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_0__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net464 (.A(clknet_0_net464),
    .X(clknet_1_1__leaf_net464));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net587 (.A(net587),
    .X(clknet_0_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_0__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_1__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net582 (.A(net582),
    .X(clknet_0_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_0__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net582 (.A(clknet_0_net582),
    .X(clknet_1_1__leaf_net582));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net695 (.A(net695),
    .X(clknet_0_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_0__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net695 (.A(clknet_0_net695),
    .X(clknet_1_1__leaf_net695));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net816 (.A(net816),
    .X(clknet_0_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net816 (.A(clknet_0_net816),
    .X(clknet_1_0__leaf_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net816 (.A(clknet_0_net816),
    .X(clknet_1_1__leaf_net816));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net333 (.A(net333),
    .X(clknet_0_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_0__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net333 (.A(clknet_0_net333),
    .X(clknet_1_1__leaf_net333));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net300 (.A(net300),
    .X(clknet_0_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_0__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net300 (.A(clknet_0_net300),
    .X(clknet_1_1__leaf_net300));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net963 (.A(net963),
    .X(clknet_0_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_1__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net869 (.A(net869),
    .X(clknet_0_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net869 (.A(clknet_0_net869),
    .X(clknet_1_0__leaf_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net869 (.A(clknet_0_net869),
    .X(clknet_1_1__leaf_net869));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net498 (.A(net498),
    .X(clknet_0_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_0__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net498 (.A(clknet_0_net498),
    .X(clknet_1_1__leaf_net498));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net314 (.A(net314),
    .X(clknet_0_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net314 (.A(clknet_0_net314),
    .X(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net287 (.A(net287),
    .X(clknet_0_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_0__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net287 (.A(clknet_0_net287),
    .X(clknet_1_1__leaf_net287));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net313 (.A(net313),
    .X(clknet_0_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_0__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net309 (.A(net309),
    .X(clknet_0_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_0__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_1__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net290 (.A(net290),
    .X(clknet_0_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net290 (.A(clknet_0_net290),
    .X(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net903 (.A(net903),
    .X(clknet_0_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net903 (.A(clknet_0_net903),
    .X(clknet_1_0__leaf_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net903 (.A(clknet_0_net903),
    .X(clknet_1_1__leaf_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net586 (.A(net586),
    .X(clknet_0_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_0__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_1__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net886 (.A(net886),
    .X(clknet_0_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_0__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_1__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net885 (.A(net885),
    .X(clknet_0_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_0__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_1__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net680 (.A(net680),
    .X(clknet_0_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_0__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net680 (.A(clknet_0_net680),
    .X(clknet_1_1__leaf_net680));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net679 (.A(net679),
    .X(clknet_0_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_0__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net679 (.A(clknet_0_net679),
    .X(clknet_1_1__leaf_net679));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net681 (.A(net681),
    .X(clknet_0_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_1__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net851 (.A(net851),
    .X(clknet_0_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net851 (.A(clknet_0_net851),
    .X(clknet_1_0__leaf_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net851 (.A(clknet_0_net851),
    .X(clknet_1_1__leaf_net851));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net850 (.A(net850),
    .X(clknet_0_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net850 (.A(clknet_0_net850),
    .X(clknet_1_0__leaf_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net850 (.A(clknet_0_net850),
    .X(clknet_1_1__leaf_net850));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net830 (.A(net830),
    .X(clknet_0_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net830 (.A(clknet_0_net830),
    .X(clknet_1_0__leaf_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net830 (.A(clknet_0_net830),
    .X(clknet_1_1__leaf_net830));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net219 (.A(net219),
    .X(clknet_0_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_0__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net219 (.A(clknet_0_net219),
    .X(clknet_1_1__leaf_net219));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net230 (.A(net230),
    .X(clknet_0_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_0__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net230 (.A(clknet_0_net230),
    .X(clknet_1_1__leaf_net230));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net218 (.A(net218),
    .X(clknet_0_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_0__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net218 (.A(clknet_0_net218),
    .X(clknet_1_1__leaf_net218));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net217 (.A(net217),
    .X(clknet_0_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_0__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net217 (.A(clknet_0_net217),
    .X(clknet_1_1__leaf_net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net216 (.A(net216),
    .X(clknet_0_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_0__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net216 (.A(clknet_0_net216),
    .X(clknet_1_1__leaf_net216));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net828 (.A(net828),
    .X(clknet_0_net828));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net828 (.A(clknet_0_net828),
    .X(clknet_1_0__leaf_net828));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net828 (.A(clknet_0_net828),
    .X(clknet_1_1__leaf_net828));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net127),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1009),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net127),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net1011),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1012),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net116),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net249),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net20),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1016),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net20),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net123),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net27),
    .X(net1020));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer13 (.A(net27),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net117),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net712),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net712),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net1024),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1024),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net982),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net6),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1028),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net947),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1030),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net947),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net42),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net1033),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1034),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net42),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net42),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net42),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net601),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net1039),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net210),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net207),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net1042),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net1042),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net14),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net848),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net916),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net847),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net70),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net203),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net838),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net807),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net417),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net223),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net422),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net351),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net846),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net652),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net346),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net414),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net827),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net875),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net225),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net209),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net598),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net883),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net824),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net788),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net796),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net732),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net837),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net338),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net353),
    .X(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_Y (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap89_A (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_RESET_B (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1_N (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1_N (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1_N (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SET_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Y (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_Y (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_Y (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_SCE (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A4 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_Y (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_Y (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_SET_B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_SCE (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCE (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_Y (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_D (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_RESET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_Y (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_SCE (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B1_N (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A3 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A4 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_Y (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_SCD (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A4 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1_N (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_D (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_Y (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_SET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCE (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_Q_N (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_SCE (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_Q (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_B1_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_RESET_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_Y (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_Y (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap60_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_D (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_Y (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_Y (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SCD (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A4 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_Y (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_Y (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A4 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_B1_N (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_SET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_SCD (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_Y (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap75_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B1_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_Y (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_B1_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A3 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_Y (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_SCD (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCE (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_SCE (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A0 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_SCD (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_SCE (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_Y (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_D (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_Y (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A3 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_SCE (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_SCD (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_SCD (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_SCD (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_D (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_RESET_B (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCD (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A4 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_SCD (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A2 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A3 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_SCE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_SCE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_S0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_Q_N (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCE (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_Q (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold67_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_S0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A4 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S0 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_SCD (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_SCD (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_X (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B1_N (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A0 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCD (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_RESET_B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_SCE (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_S0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCD (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1_N (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_Y (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_SCD (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_SCE (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_Y (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_D (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q_N (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCD (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_Q (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_RESET_B (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_SCE (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_Q (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_Q_N (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1_N (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_Q (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_X (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_Y (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_RESET_B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_Q (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_RESET_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_X (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A3 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_SCD (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_B1_N (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_Y (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_SET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Y (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_S1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCD (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_B1_N (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A4 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1_N (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A0 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B1_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_B1_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SCD (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A0 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A2 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_Y (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_X (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_SCE (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_RESET_B (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SCD (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SCD (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A4 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_X (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_SET_B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SCE (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_X (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_X (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_RESET_B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A3 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A4 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_Y (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_D (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A4 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_X (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SCD (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_X (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A3 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_RESET_B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_D (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_X (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_X (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S0 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_SET_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SCE (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_SCE (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_RESET_B (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_X (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_Y (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B1_N (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A4 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_Q (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_SET_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_B1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_Q (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_SET_B (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q_N (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A4 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1_N (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_Q (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q_N (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_S1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_B1_N (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A3 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_Q (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_Q (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_Q (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B1_N (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_Q (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_Q_N (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_Q (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_Q (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_SET_B (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B1_N (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_Y (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A4 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_B1_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B1_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B1_N (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_B1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_B1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_Q (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_SCD (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_SCD (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B1_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_S0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B1_N (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A4 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B1_N (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_B1 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_A2 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A1 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_B1_N (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B1_N (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A1 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_RESET_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_Q (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_S1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_Y (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_B1_N (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_SCD (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_Q (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_B1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_Q (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_RESET_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_RESET_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_SET_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_SCD (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_SCE (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_Q (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap66_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_S0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A4 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_Y (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A4 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B1_N (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_Y (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_Q (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_Q (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap68_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_Y (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_Q (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_SET_B (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A2 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap61_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_SET_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_Y (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A3 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCE (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A4 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCE (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_RESET_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_B1_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_SCE (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_S1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_SCD (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B1_N (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B1_N (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_SCE (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_D (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap60_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap59_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SET_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap61_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A2 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_B1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire63_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SET_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A4 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A4 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_SCE (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_B1_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap66_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SCD (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap68_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1_N (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1_N (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B1_N (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SET_B (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCE (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap73_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SET_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_RESET_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_SCE (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap75_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap76_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A4 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B1_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_SET_B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_SCD (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_SCD (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCD (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_SCD (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A4 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SET_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_RESET_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A4 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_S0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_SCD (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_SCD (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A3 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap87_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_D (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap89_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s885_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_SLEEP_B (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s874_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s875_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s877_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s882_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s846_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A1 (.DIODE(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net408_X (.DIODE(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net964_A (.DIODE(clknet_0_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net964_A (.DIODE(clknet_0_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net964_X (.DIODE(clknet_0_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_B1_N (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1_N (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_SET_B (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_SET_B (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SET_B (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B1 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A2 (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net964_X (.DIODE(clknet_1_0__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_S0 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A1 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B1 (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net964_X (.DIODE(clknet_1_1__leaf_net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCE (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S0 (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net304_X (.DIODE(clknet_1_0__leaf_net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SCE (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net315_X (.DIODE(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A4 (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_S1 (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A2 (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A0 (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net315_X (.DIODE(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A4 (.DIODE(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_B1 (.DIODE(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_S1 (.DIODE(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net314_X (.DIODE(clknet_1_0__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCD (.DIODE(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net314_X (.DIODE(clknet_1_1__leaf_net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_SET_B (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A0 (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_B1 (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net290_X (.DIODE(clknet_1_0__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A4 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A3 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_S0 (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net290_X (.DIODE(clknet_1_1__leaf_net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_X (.DIODE(net1019));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net515),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net515),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net515),
    .X(net1078));
 sky130_fd_sc_hd__xnor2_1 clone43 (.A(net925),
    .B(net921),
    .Y(net1079));
 sky130_fd_sc_hd__xnor2_1 clone44 (.A(net509),
    .B(net508),
    .Y(net1080));
 sky130_fd_sc_hd__a21bo_1 clone45 (.A1(net112),
    .A2(net120),
    .B1_N(net121),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_1 clone46 (.A(net990),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net33),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net33),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net151),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net1085),
    .X(net1086));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
