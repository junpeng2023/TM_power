module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net644;
 wire clknet_1_0__leaf_net644;
 wire clknet_1_1__leaf_net644;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net660;
 wire clknet_1_0__leaf_net660;
 wire clknet_1_1__leaf_net660;
 wire clknet_0_net661;
 wire clknet_1_0__leaf_net661;
 wire clknet_1_1__leaf_net661;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net653;
 wire clknet_1_0__leaf_net653;
 wire clknet_1_1__leaf_net653;
 wire clknet_0_net590;
 wire clknet_1_0__leaf_net590;
 wire clknet_1_1__leaf_net590;
 wire clknet_0_net751;
 wire clknet_1_0__leaf_net751;
 wire clknet_1_1__leaf_net751;
 wire clknet_0_net594;
 wire clknet_1_0__leaf_net594;
 wire clknet_1_1__leaf_net594;
 wire clknet_0_net587;
 wire clknet_1_0__leaf_net587;
 wire clknet_1_1__leaf_net587;
 wire clknet_0_net743;
 wire clknet_1_0__leaf_net743;
 wire clknet_1_1__leaf_net743;
 wire clknet_0_net689;
 wire clknet_1_0__leaf_net689;
 wire clknet_1_1__leaf_net689;
 wire clknet_0_net589;
 wire clknet_1_0__leaf_net589;
 wire clknet_1_1__leaf_net589;
 wire clknet_0_net564;
 wire clknet_1_0__leaf_net564;
 wire clknet_1_1__leaf_net564;
 wire clknet_0_net577;
 wire clknet_1_0__leaf_net577;
 wire clknet_1_1__leaf_net577;
 wire clknet_0_net668;
 wire clknet_1_0__leaf_net668;
 wire clknet_1_1__leaf_net668;
 wire clknet_0_net571;
 wire clknet_1_0__leaf_net571;
 wire clknet_1_1__leaf_net571;
 wire clknet_0_net575;
 wire clknet_1_0__leaf_net575;
 wire clknet_1_1__leaf_net575;
 wire clknet_0_net670;
 wire clknet_1_0__leaf_net670;
 wire clknet_1_1__leaf_net670;
 wire clknet_0_net678;
 wire clknet_1_0__leaf_net678;
 wire clknet_1_1__leaf_net678;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net586;
 wire clknet_1_0__leaf_net586;
 wire clknet_1_1__leaf_net586;
 wire clknet_0_net584;
 wire clknet_1_0__leaf_net584;
 wire clknet_1_1__leaf_net584;
 wire clknet_0_net583;
 wire clknet_1_0__leaf_net583;
 wire clknet_1_1__leaf_net583;
 wire clknet_0_net565;
 wire clknet_1_0__leaf_net565;
 wire clknet_1_1__leaf_net565;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net542;
 wire clknet_1_0__leaf_net542;
 wire clknet_1_1__leaf_net542;
 wire clknet_0_net649;
 wire clknet_1_0__leaf_net649;
 wire clknet_1_1__leaf_net649;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net549;
 wire clknet_1_0__leaf_net549;
 wire clknet_1_1__leaf_net549;
 wire clknet_0_net555;
 wire clknet_1_0__leaf_net555;
 wire clknet_1_1__leaf_net555;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net556;
 wire clknet_1_0__leaf_net556;
 wire clknet_1_1__leaf_net556;
 wire clknet_0_net551;
 wire clknet_1_0__leaf_net551;
 wire clknet_1_1__leaf_net551;
 wire clknet_0_net548;
 wire clknet_1_0__leaf_net548;
 wire clknet_1_1__leaf_net548;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net547;
 wire clknet_1_0__leaf_net547;
 wire clknet_1_1__leaf_net547;
 wire clknet_0_net545;
 wire clknet_1_0__leaf_net545;
 wire clknet_1_1__leaf_net545;
 wire clknet_0_net335;
 wire clknet_1_0__leaf_net335;
 wire clknet_1_1__leaf_net335;
 wire clknet_0_net336;
 wire clknet_1_0__leaf_net336;
 wire clknet_1_1__leaf_net336;
 wire clknet_0_net347;
 wire clknet_1_0__leaf_net347;
 wire clknet_1_1__leaf_net347;
 wire clknet_0_net338;
 wire clknet_1_0__leaf_net338;
 wire clknet_1_1__leaf_net338;
 wire clknet_0_net337;
 wire clknet_1_0__leaf_net337;
 wire clknet_1_1__leaf_net337;
 wire clknet_0_net334;
 wire clknet_1_0__leaf_net334;
 wire clknet_1_1__leaf_net334;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;

 sky130_fd_sc_hd__and3_1 c100 (.A(net73),
    .B(net72),
    .C(net74),
    .X(net77));
 sky130_fd_sc_hd__and3_1 c101 (.A(net61),
    .B(net74),
    .C(net72),
    .X(net78));
 sky130_fd_sc_hd__and3_1 c102 (.A(net78),
    .B(net76),
    .C(net74),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net77),
    .A1(net72),
    .A2(net71),
    .A3(net68),
    .S0(net63),
    .S1(net755),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net69),
    .A1(net79),
    .A2(net76),
    .A3(net63),
    .S0(net755),
    .S1(net705),
    .X(net81));
 sky130_fd_sc_hd__buf_1 c105 (.A(net706),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 c106 (.A(net55),
    .X(net83));
 sky130_fd_sc_hd__and2_1 c107 (.A(net82),
    .B(net83),
    .X(net84));
 sky130_fd_sc_hd__and2_0 c108 (.A(net84),
    .B(net83),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 c109 (.A(net83),
    .X(net86));
 sky130_fd_sc_hd__and2_0 c110 (.A(net85),
    .B(net83),
    .X(net87));
 sky130_fd_sc_hd__and2_1 c111 (.A(net86),
    .B(net84),
    .X(net88));
 sky130_fd_sc_hd__and2_0 c112 (.A(net82),
    .B(net88),
    .X(net89));
 sky130_fd_sc_hd__and2_0 c113 (.A(net83),
    .B(net88),
    .X(net90));
 sky130_fd_sc_hd__and2_1 c114 (.A(net84),
    .B(net82),
    .X(net91));
 sky130_fd_sc_hd__and3_1 c115 (.A(net88),
    .B(net91),
    .C(net83),
    .X(net92));
 sky130_fd_sc_hd__and2_1 c116 (.A(net89),
    .B(net91),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c117 (.A(net93),
    .B(net88),
    .X(net94));
 sky130_fd_sc_hd__and3_1 c118 (.A(net92),
    .B(net82),
    .C(net93),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 c119 (.A0(net90),
    .A1(net93),
    .A2(net84),
    .A3(net95),
    .S0(net92),
    .S1(net94),
    .X(net96));
 sky130_fd_sc_hd__and3_1 c120 (.A(net94),
    .B(net91),
    .C(net93),
    .X(net97));
 sky130_fd_sc_hd__and3_1 c121 (.A(net91),
    .B(net93),
    .C(net95),
    .X(net98));
 sky130_fd_sc_hd__and3_1 c122 (.A(net87),
    .B(net98),
    .C(net96),
    .X(net99));
 sky130_fd_sc_hd__and3_1 c123 (.A(net97),
    .B(net95),
    .C(net96),
    .X(net100));
 sky130_fd_sc_hd__and2_0 c124 (.A(net96),
    .B(net99),
    .X(net101));
 sky130_fd_sc_hd__or4bb_1 c125 (.A(net101),
    .B(net100),
    .C_N(net95),
    .D_N(net82),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 c126 (.A(in0),
    .X(net103));
 sky130_fd_sc_hd__and2_0 c127 (.A(net103),
    .B(net735),
    .X(net104));
 sky130_fd_sc_hd__and2_0 c128 (.A(net104),
    .B(net103),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 c129 (.A(in12),
    .X(net106));
 sky130_fd_sc_hd__and2_0 c130 (.A(net106),
    .B(net734),
    .X(net107));
 sky130_fd_sc_hd__and2_0 c131 (.A(net722),
    .B(net726),
    .X(net108));
 sky130_fd_sc_hd__and2_0 c132 (.A(net107),
    .B(net720),
    .X(net109));
 sky130_fd_sc_hd__and2_0 c133 (.A(net733),
    .B(net108),
    .X(net110));
 sky130_fd_sc_hd__and2_1 c134 (.A(net110),
    .B(net105),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c135 (.A(net106),
    .B(net111),
    .C(net104),
    .X(net112));
 sky130_fd_sc_hd__and3_1 c136 (.A(net108),
    .B(net721),
    .C(net111),
    .X(net113));
 sky130_fd_sc_hd__and3_1 c137 (.A(net105),
    .B(net110),
    .C(net111),
    .X(net114));
 sky130_fd_sc_hd__and2_0 c138 (.A(net111),
    .B(net114),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c139 (.A(net113),
    .B(net112),
    .C(net109),
    .X(net116));
 sky130_fd_sc_hd__and3_1 c140 (.A(net116),
    .B(net111),
    .C(net109),
    .X(net117));
 sky130_fd_sc_hd__and3_1 c141 (.A(net114),
    .B(net113),
    .C(net111),
    .X(net118));
 sky130_fd_sc_hd__or4bb_1 c142 (.A(net112),
    .B(net717),
    .C_N(net116),
    .D_N(net117),
    .X(net119));
 sky130_fd_sc_hd__and3_1 c143 (.A(net115),
    .B(net118),
    .C(net119),
    .X(net120));
 sky130_fd_sc_hd__and3_1 c144 (.A(net109),
    .B(net119),
    .C(net113),
    .X(net121));
 sky130_fd_sc_hd__a2111o_1 c145 (.A1(net120),
    .A2(net738),
    .B1(net121),
    .C1(net111),
    .D1(net117),
    .X(net122));
 sky130_fd_sc_hd__and3_1 c146 (.A(net121),
    .B(net122),
    .C(net111),
    .X(net123));
 sky130_fd_sc_hd__buf_1 c147 (.A(net7),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 c148 (.A(net124),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 c149 (.A(net125),
    .X(net126));
 sky130_fd_sc_hd__and2_2 c150 (.A(net16),
    .B(net125),
    .X(net127));
 sky130_fd_sc_hd__and2_0 c151 (.A(net127),
    .B(net125),
    .X(net128));
 sky130_fd_sc_hd__and2_0 c152 (.A(net124),
    .B(net127),
    .X(net129));
 sky130_fd_sc_hd__and2_0 c153 (.A(net127),
    .B(net125),
    .X(net130));
 sky130_fd_sc_hd__and3_1 c154 (.A(net128),
    .B(net124),
    .C(net127),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c155 (.A(net125),
    .B(net131),
    .X(net132));
 sky130_fd_sc_hd__and2_0 c156 (.A(net132),
    .B(net131),
    .X(net133));
 sky130_fd_sc_hd__and3_1 c157 (.A(net2),
    .B(net127),
    .C(net131),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c158 (.A0(net131),
    .A1(net127),
    .A2(net123),
    .A3(net134),
    .S0(net125),
    .S1(net132),
    .X(net135));
 sky130_fd_sc_hd__and2_0 c159 (.A(net130),
    .B(net132),
    .X(net136));
 sky130_fd_sc_hd__and2_0 c160 (.A(net134),
    .B(net124),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c161 (.A0(net136),
    .A1(net134),
    .A2(net127),
    .A3(net132),
    .S0(net131),
    .S1(net125),
    .X(net138));
 sky130_fd_sc_hd__and3_1 c162 (.A(net129),
    .B(net124),
    .C(net134),
    .X(net139));
 sky130_fd_sc_hd__or4bb_1 c163 (.A(net125),
    .B(net139),
    .C_N(net134),
    .D_N(net123),
    .X(net140));
 sky130_fd_sc_hd__and2_0 c164 (.A(net138),
    .B(net139),
    .X(net141));
 sky130_fd_sc_hd__a2111o_1 c165 (.A1(net137),
    .A2(net141),
    .B1(net139),
    .C1(net127),
    .D1(net131),
    .X(net142));
 sky130_fd_sc_hd__and3_1 c166 (.A(net126),
    .B(net142),
    .C(net117),
    .X(net143));
 sky130_fd_sc_hd__a2111o_1 c167 (.A1(net143),
    .A2(net135),
    .B1(net139),
    .C1(net125),
    .D1(net127),
    .X(net144));
 sky130_fd_sc_hd__buf_1 c168 (.A(net26),
    .X(net145));
 sky130_fd_sc_hd__and2_0 c169 (.A(net144),
    .B(net145),
    .X(net146));
 sky130_fd_sc_hd__buf_1 c170 (.A(net145),
    .X(net147));
 sky130_fd_sc_hd__buf_1 c171 (.A(net147),
    .X(net148));
 sky130_fd_sc_hd__and2_0 c172 (.A(net148),
    .B(net147),
    .X(net149));
 sky130_fd_sc_hd__and2_0 c173 (.A(net145),
    .B(net148),
    .X(net150));
 sky130_fd_sc_hd__and2_0 c174 (.A(net148),
    .B(net149),
    .X(net151));
 sky130_fd_sc_hd__and2_0 c175 (.A(net150),
    .B(net148),
    .X(net152));
 sky130_fd_sc_hd__dfrtp_1 c176 (.CLK(clknet_4_1_0_clk),
    .D(net146),
    .RESET_B(net37),
    .Q(net153));
 sky130_fd_sc_hd__and2_1 c177 (.A(net795),
    .B(net34),
    .X(net154));
 sky130_fd_sc_hd__and2_0 c178 (.A(net145),
    .B(net154),
    .X(net155));
 sky130_fd_sc_hd__and2_0 c179 (.A(net152),
    .B(net147),
    .X(net156));
 sky130_fd_sc_hd__and2_1 c180 (.A(net149),
    .B(net154),
    .X(net157));
 sky130_fd_sc_hd__and2_0 c181 (.A(net795),
    .B(net157),
    .X(net158));
 sky130_fd_sc_hd__and2_0 c182 (.A(net151),
    .B(net157),
    .X(net159));
 sky130_fd_sc_hd__sdfbbn_1 c183 (.CLK_N(clknet_4_1_0_clk),
    .D(net155),
    .RESET_B(net159),
    .SCD(net156),
    .SCE(net154),
    .SET_B(net37),
    .Q(net161),
    .Q_N(net160));
 sky130_fd_sc_hd__and3_1 c184 (.A(net147),
    .B(net160),
    .C(net157),
    .X(net162));
 sky130_fd_sc_hd__dfrtp_1 c185 (.CLK(clknet_4_0_0_clk),
    .D(net157),
    .RESET_B(net162),
    .Q(net163));
 sky130_fd_sc_hd__dfsbp_1 c186 (.CLK(clknet_4_0_0_clk),
    .D(net154),
    .SET_B(net159),
    .Q(net165),
    .Q_N(net164));
 sky130_fd_sc_hd__dfbbn_1 c187 (.CLK_N(clknet_4_0_0_clk),
    .D(net165),
    .RESET_B(net163),
    .SET_B(net162),
    .Q(net166));
 sky130_fd_sc_hd__and3_1 c188 (.A(net163),
    .B(net166),
    .C(net164),
    .X(net167));
 sky130_fd_sc_hd__dfsbp_1 c189 (.CLK(clknet_4_0_0_clk),
    .D(net158),
    .SET_B(net60),
    .Q(net169),
    .Q_N(net168));
 sky130_fd_sc_hd__clkbuf_2 c190 (.A(net168),
    .X(net170));
 sky130_fd_sc_hd__and2_0 c191 (.A(net167),
    .B(net170),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 c192 (.A(net170),
    .X(net172));
 sky130_fd_sc_hd__and2_0 c193 (.A(net169),
    .B(net170),
    .X(net173));
 sky130_fd_sc_hd__and2_0 c194 (.A(net171),
    .B(net170),
    .X(net174));
 sky130_fd_sc_hd__and2_0 c195 (.A(net174),
    .B(net170),
    .X(net175));
 sky130_fd_sc_hd__and2_1 c196 (.A(net174),
    .B(net170),
    .X(net176));
 sky130_fd_sc_hd__and2_0 c197 (.A(net175),
    .B(net170),
    .X(net177));
 sky130_fd_sc_hd__and2_0 c198 (.A(net173),
    .B(net55),
    .X(net178));
 sky130_fd_sc_hd__and2_1 c199 (.A(net170),
    .B(net175),
    .X(net179));
 sky130_fd_sc_hd__and2_0 c200 (.A(net172),
    .B(net60),
    .X(net180));
 sky130_fd_sc_hd__and2_0 c201 (.A(net171),
    .B(net180),
    .X(net181));
 sky130_fd_sc_hd__and2_0 c202 (.A(net180),
    .B(net60),
    .X(net182));
 sky130_fd_sc_hd__and2_0 c203 (.A(net181),
    .B(net182),
    .X(net183));
 sky130_fd_sc_hd__and2_0 c204 (.A(net177),
    .B(net183),
    .X(net184));
 sky130_fd_sc_hd__and2_0 c205 (.A(net182),
    .B(net177),
    .X(net185));
 sky130_fd_sc_hd__and2_0 c206 (.A(net172),
    .B(net185),
    .X(net186));
 sky130_fd_sc_hd__and2_1 c207 (.A(net184),
    .B(net179),
    .X(net187));
 sky130_fd_sc_hd__a2111o_1 c208 (.A1(net185),
    .A2(net186),
    .B1(net187),
    .C1(net44),
    .D1(net170),
    .X(net188));
 sky130_fd_sc_hd__and2_0 c209 (.A(net178),
    .B(net188),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 c210 (.A(net189),
    .X(net190));
 sky130_fd_sc_hd__and2_2 c211 (.A(net187),
    .B(net755),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 c212 (.A(net191),
    .X(net192));
 sky130_fd_sc_hd__and2_1 c213 (.A(net190),
    .B(net191),
    .X(net193));
 sky130_fd_sc_hd__and2_0 c214 (.A(net192),
    .B(net190),
    .X(net194));
 sky130_fd_sc_hd__dfstp_1 c215 (.CLK(clknet_4_2_0_clk),
    .D(net193),
    .SET_B(net191),
    .Q(net195));
 sky130_fd_sc_hd__and2_0 c216 (.A(net191),
    .B(net195),
    .X(net196));
 sky130_fd_sc_hd__dfstp_1 c217 (.CLK(clknet_4_2_0_clk),
    .D(net194),
    .SET_B(net191),
    .Q(net197));
 sky130_fd_sc_hd__and2_0 c218 (.A(net75),
    .B(net192),
    .X(net198));
 sky130_fd_sc_hd__dfbbn_1 c219 (.CLK_N(clknet_4_2_0_clk),
    .D(net183),
    .RESET_B(net193),
    .SET_B(net755),
    .Q(net200),
    .Q_N(net199));
 sky130_fd_sc_hd__and2_0 c220 (.A(net197),
    .B(net200),
    .X(net201));
 sky130_fd_sc_hd__and2_0 c221 (.A(net196),
    .B(net200),
    .X(net202));
 sky130_fd_sc_hd__and2_1 c222 (.A(net755),
    .B(net200),
    .X(net203));
 sky130_fd_sc_hd__sdfbbn_1 c223 (.CLK_N(clknet_4_2_0_clk),
    .D(net201),
    .RESET_B(net194),
    .SCD(net191),
    .SCE(net199),
    .SET_B(net203),
    .Q(net204));
 sky130_fd_sc_hd__and2_1 c224 (.A(net204),
    .B(net203),
    .X(net205));
 sky130_fd_sc_hd__dfstp_1 c225 (.CLK(clknet_4_8_0_clk),
    .D(net198),
    .SET_B(net205),
    .Q(net206));
 sky130_fd_sc_hd__or4bb_1 c226 (.A(net202),
    .B(net205),
    .C_N(net196),
    .D_N(net176),
    .X(net207));
 sky130_fd_sc_hd__dfbbp_1 c227 (.CLK(clknet_4_8_0_clk),
    .D(net207),
    .RESET_B(net205),
    .SET_B(net202),
    .Q(net209),
    .Q_N(net208));
 sky130_fd_sc_hd__sdfbbp_1 c228 (.CLK(clknet_4_2_0_clk),
    .D(net195),
    .RESET_B(net209),
    .SCD(net193),
    .SCE(net199),
    .SET_B(net191),
    .Q(net211),
    .Q_N(net210));
 sky130_fd_sc_hd__a2111o_1 c229 (.A1(net179),
    .A2(net211),
    .B1(net209),
    .C1(net199),
    .D1(net67),
    .X(net212));
 sky130_fd_sc_hd__sdfbbn_1 c230 (.CLK_N(clknet_4_8_0_clk),
    .D(net212),
    .RESET_B(net195),
    .SCD(net207),
    .SCE(net210),
    .SET_B(net208),
    .Q(net214),
    .Q_N(net213));
 sky130_fd_sc_hd__clkbuf_1 c231 (.A(net206),
    .X(net215));
 sky130_fd_sc_hd__dlymetal6s2s_1 c232 (.A(net102),
    .X(net216));
 sky130_fd_sc_hd__dlrbn_1 c233 (.D(net215),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net216),
    .Q(net753),
    .Q_N(net217));
 sky130_fd_sc_hd__and2_0 c234 (.A(net215),
    .B(net217),
    .X(net218));
 sky130_fd_sc_hd__and2_0 c235 (.A(net215),
    .B(net213),
    .X(net219));
 sky130_fd_sc_hd__dlrbn_1 c236 (.D(net216),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net217),
    .Q(net220));
 sky130_fd_sc_hd__dlrbp_1 c237 (.D(net220),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net216),
    .Q(net222),
    .Q_N(net221));
 sky130_fd_sc_hd__and2_0 c238 (.A(net218),
    .B(net222),
    .X(net223));
 sky130_fd_sc_hd__sdfxbp_1 c239 (.CLK(clknet_4_8_0_clk),
    .D(net787),
    .SCD(net216),
    .SCE(net217),
    .Q(net225),
    .Q_N(net224));
 sky130_fd_sc_hd__and3_1 c240 (.A(net223),
    .B(net225),
    .C(net221),
    .X(net226));
 sky130_fd_sc_hd__dlrbp_1 c241 (.D(net216),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net222),
    .Q(net227));
 sky130_fd_sc_hd__and2_0 c242 (.A(net222),
    .B(net753),
    .X(net228));
 sky130_fd_sc_hd__and2_0 c243 (.A(net226),
    .B(net224),
    .X(net229));
 sky130_fd_sc_hd__sdfxbp_1 c244 (.CLK(clknet_4_8_0_clk),
    .D(net228),
    .SCD(net216),
    .SCE(net753),
    .Q(net231),
    .Q_N(net230));
 sky130_fd_sc_hd__and2_0 c245 (.A(net229),
    .B(net224),
    .X(net232));
 sky130_fd_sc_hd__and3_1 c246 (.A(net231),
    .B(net753),
    .C(net223),
    .X(net233));
 sky130_fd_sc_hd__and3_1 c247 (.A(net233),
    .B(net225),
    .C(net221),
    .X(net234));
 sky130_fd_sc_hd__and3_1 c248 (.A(net227),
    .B(net234),
    .C(net224),
    .X(net235));
 sky130_fd_sc_hd__and3_1 c249 (.A(net234),
    .B(net235),
    .C(net230),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c25 (.A(net731),
    .B(net739),
    .X(net0));
 sky130_fd_sc_hd__and3_1 c250 (.A(net225),
    .B(net235),
    .C(net234),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net237),
    .A1(net231),
    .A2(net214),
    .A3(net235),
    .S0(net217),
    .S1(net221),
    .X(net238));
 sky130_fd_sc_hd__buf_1 c252 (.A(net117),
    .X(net239));
 sky130_fd_sc_hd__buf_1 c253 (.A(net239),
    .X(net240));
 sky130_fd_sc_hd__buf_1 c254 (.A(net239),
    .X(net241));
 sky130_fd_sc_hd__and2_0 c255 (.A(net240),
    .B(net123),
    .X(net242));
 sky130_fd_sc_hd__and2_0 c256 (.A(net239),
    .B(net241),
    .X(net243));
 sky130_fd_sc_hd__and2_1 c257 (.A(net240),
    .B(net241),
    .X(net244));
 sky130_fd_sc_hd__and2_1 c258 (.A(net241),
    .B(net724),
    .X(net245));
 sky130_fd_sc_hd__and2_0 c259 (.A(net245),
    .B(net243),
    .X(net246));
 sky130_fd_sc_hd__and2_0 c26 (.A(net729),
    .B(net727),
    .X(net1));
 sky130_fd_sc_hd__and2_0 c260 (.A(net241),
    .B(net240),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c261 (.A(net246),
    .B(net239),
    .C(net247),
    .X(net248));
 sky130_fd_sc_hd__and2_0 c262 (.A(net245),
    .B(net247),
    .X(net249));
 sky130_fd_sc_hd__and3_2 c263 (.A(net247),
    .B(net244),
    .C(net245),
    .X(net250));
 sky130_fd_sc_hd__or4bb_1 c264 (.A(net242),
    .B(net241),
    .C_N(net244),
    .D_N(net245),
    .X(net251));
 sky130_fd_sc_hd__and2_0 c265 (.A(net117),
    .B(net250),
    .X(net252));
 sky130_fd_sc_hd__or4bb_1 c266 (.A(net243),
    .B(net249),
    .C_N(net252),
    .D_N(net250),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c267 (.A0(net244),
    .A1(net240),
    .A2(net246),
    .A3(net123),
    .S0(net241),
    .S1(net250),
    .X(net254));
 sky130_fd_sc_hd__and2_0 c268 (.A(net246),
    .B(net250),
    .X(net255));
 sky130_fd_sc_hd__and3_1 c269 (.A(net254),
    .B(net255),
    .C(net250),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c27 (.A(net731),
    .B(net719),
    .C(net730),
    .X(net2));
 sky130_fd_sc_hd__or4bb_1 c270 (.A(net252),
    .B(net256),
    .C_N(net253),
    .D_N(net250),
    .X(net257));
 sky130_fd_sc_hd__or4bb_1 c271 (.A(net253),
    .B(net251),
    .C_N(net256),
    .D_N(net244),
    .X(net258));
 sky130_fd_sc_hd__or4bb_1 c272 (.A(net258),
    .B(net257),
    .C_N(net251),
    .D_N(net256),
    .X(net259));
 sky130_fd_sc_hd__buf_1 c273 (.A(net123),
    .X(net260));
 sky130_fd_sc_hd__and2_1 c274 (.A(net260),
    .B(net250),
    .X(net261));
 sky130_fd_sc_hd__and2_0 c275 (.A(net260),
    .B(net261),
    .X(net262));
 sky130_fd_sc_hd__and2_1 c276 (.A(net262),
    .B(net261),
    .X(net263));
 sky130_fd_sc_hd__and2_0 c277 (.A(net133),
    .B(net261),
    .X(net264));
 sky130_fd_sc_hd__and3_1 c278 (.A(net123),
    .B(net260),
    .C(net261),
    .X(net265));
 sky130_fd_sc_hd__and2_1 c279 (.A(net263),
    .B(net265),
    .X(net266));
 sky130_fd_sc_hd__and3_1 c28 (.A(net1),
    .B(net728),
    .C(net730),
    .X(net3));
 sky130_fd_sc_hd__and2_0 c280 (.A(net140),
    .B(net261),
    .X(net267));
 sky130_fd_sc_hd__and2_1 c281 (.A(net267),
    .B(net262),
    .X(net268));
 sky130_fd_sc_hd__and2_0 c282 (.A(net268),
    .B(net265),
    .X(net269));
 sky130_fd_sc_hd__and3_1 c283 (.A(net260),
    .B(net265),
    .C(net263),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c284 (.A(net265),
    .B(net264),
    .C(net268),
    .X(net271));
 sky130_fd_sc_hd__or4bb_2 c285 (.A(net264),
    .B(net271),
    .C_N(net270),
    .D_N(net263),
    .X(net272));
 sky130_fd_sc_hd__and2_1 c286 (.A(net269),
    .B(net263),
    .X(net273));
 sky130_fd_sc_hd__and3_1 c287 (.A(net271),
    .B(net273),
    .C(net268),
    .X(net274));
 sky130_fd_sc_hd__and2_1 c288 (.A(net273),
    .B(net271),
    .X(net275));
 sky130_fd_sc_hd__a2111o_1 c289 (.A1(net274),
    .A2(net271),
    .B1(net263),
    .C1(net272),
    .D1(net260),
    .X(net276));
 sky130_fd_sc_hd__and2_0 c29 (.A(net730),
    .B(net0),
    .X(net4));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net270),
    .A1(net272),
    .A2(net276),
    .A3(net273),
    .S0(net271),
    .S1(net259),
    .X(net277));
 sky130_fd_sc_hd__and3_1 c291 (.A(net261),
    .B(net273),
    .C(net707),
    .X(net278));
 sky130_fd_sc_hd__and3_1 c292 (.A(net278),
    .B(net268),
    .C(net273),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net276),
    .A1(net275),
    .A2(net261),
    .A3(net270),
    .S0(net279),
    .S1(net707),
    .X(net280));
 sky130_fd_sc_hd__buf_1 c294 (.A(net156),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 c295 (.A(net34),
    .X(net282));
 sky130_fd_sc_hd__buf_1 c296 (.A(net272),
    .X(net283));
 sky130_fd_sc_hd__dlrtn_1 c297 (.D(net279),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net283),
    .Q(net284));
 sky130_fd_sc_hd__and2_1 c298 (.A(net284),
    .B(net281),
    .X(net285));
 sky130_fd_sc_hd__and2_1 c299 (.A(net281),
    .B(net283),
    .X(net286));
 sky130_fd_sc_hd__and2_1 c30 (.A(net732),
    .B(net723),
    .X(net5));
 sky130_fd_sc_hd__dlrtn_1 c300 (.D(net284),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net286),
    .Q(net287));
 sky130_fd_sc_hd__sdfxtp_1 c301 (.CLK(clknet_4_4_0_clk),
    .D(net287),
    .SCD(net286),
    .SCE(net283),
    .Q(net288));
 sky130_fd_sc_hd__and3_1 c302 (.A(net282),
    .B(net288),
    .C(net285),
    .X(net289));
 sky130_fd_sc_hd__and3_1 c303 (.A(net289),
    .B(net281),
    .C(net288),
    .X(net290));
 sky130_fd_sc_hd__and3_1 c304 (.A(net281),
    .B(net285),
    .C(net284),
    .X(net291));
 sky130_fd_sc_hd__sdfxtp_1 c305 (.CLK(clknet_4_4_0_clk),
    .D(net285),
    .SCD(net286),
    .SCE(net291),
    .Q(net292));
 sky130_fd_sc_hd__and3_1 c306 (.A(net803),
    .B(net288),
    .C(net291),
    .X(net293));
 sky130_fd_sc_hd__and3_1 c307 (.A(net161),
    .B(net291),
    .C(net285),
    .X(net294));
 sky130_fd_sc_hd__sdfxtp_1 c308 (.CLK(clknet_4_1_0_clk),
    .D(net290),
    .SCD(net293),
    .SCE(net284),
    .Q(net295));
 sky130_fd_sc_hd__a2111o_1 c309 (.A1(net295),
    .A2(net291),
    .B1(net281),
    .C1(net288),
    .D1(net800),
    .X(net296));
 sky130_fd_sc_hd__and2_0 c31 (.A(net8),
    .B(net2),
    .X(net6));
 sky130_fd_sc_hd__dfbbn_1 c310 (.CLK_N(clknet_4_1_0_clk),
    .D(net283),
    .RESET_B(net286),
    .SET_B(net288),
    .Q(net298),
    .Q_N(net297));
 sky130_fd_sc_hd__dfbbn_1 c311 (.CLK_N(clknet_4_1_0_clk),
    .D(net778),
    .RESET_B(net296),
    .SET_B(net290),
    .Q(net299));
 sky130_fd_sc_hd__and3_1 c312 (.A(net288),
    .B(net285),
    .C(net297),
    .X(net300));
 sky130_fd_sc_hd__and3_1 c313 (.A(net299),
    .B(net283),
    .C(net34),
    .X(net301));
 sky130_fd_sc_hd__dfbbp_1 c314 (.CLK(clknet_4_1_0_clk),
    .D(net300),
    .RESET_B(net294),
    .SET_B(net301),
    .Q(net303),
    .Q_N(net302));
 sky130_fd_sc_hd__dlymetal6s2s_1 c315 (.A(net189),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 c316 (.A(net304),
    .X(net305));
 sky130_fd_sc_hd__and2_2 c317 (.A(net44),
    .B(net304),
    .X(net306));
 sky130_fd_sc_hd__dlrtn_1 c318 (.D(net304),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net305),
    .Q(net307));
 sky130_fd_sc_hd__dlrtp_1 c319 (.D(net305),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net306),
    .Q(net308));
 sky130_fd_sc_hd__a2111o_2 c32 (.A1(net3),
    .A2(net5),
    .B1(net4),
    .C1(net730),
    .D1(net732),
    .X(net7));
 sky130_fd_sc_hd__dlrtp_1 c320 (.D(net307),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net306),
    .Q(net309));
 sky130_fd_sc_hd__sdfxbp_1 c321 (.CLK(clknet_4_3_0_clk),
    .D(net304),
    .SCD(net187),
    .SCE(net306),
    .Q(net310));
 sky130_fd_sc_hd__and2_0 c322 (.A(net808),
    .B(net307),
    .X(net311));
 sky130_fd_sc_hd__dlrtp_1 c323 (.D(net301),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net304),
    .Q(net312));
 sky130_fd_sc_hd__edfxbp_1 c324 (.CLK(clknet_4_3_0_clk),
    .D(net305),
    .DE(net306),
    .Q(net313));
 sky130_fd_sc_hd__edfxtp_1 c325 (.CLK(clknet_4_2_0_clk),
    .D(net307),
    .DE(net305),
    .Q(net314));
 sky130_fd_sc_hd__sdfxbp_1 c326 (.CLK(clknet_4_3_0_clk),
    .D(net772),
    .SCD(net307),
    .SCE(net306),
    .Q(net316),
    .Q_N(net315));
 sky130_fd_sc_hd__sdfxtp_1 c327 (.CLK(clknet_4_2_0_clk),
    .D(net306),
    .SCD(net304),
    .SCE(net790),
    .Q(net317));
 sky130_fd_sc_hd__and3_1 c328 (.A(net314),
    .B(net317),
    .C(net176),
    .X(net318));
 sky130_fd_sc_hd__sdfxtp_1 c329 (.CLK(clknet_4_2_0_clk),
    .D(net780),
    .SCD(net792),
    .SCE(net305),
    .Q(net319));
 sky130_fd_sc_hd__and2_0 c33 (.A(net736),
    .B(net737),
    .X(net8));
 sky130_fd_sc_hd__and3_1 c330 (.A(net318),
    .B(net314),
    .C(net316),
    .X(net320));
 sky130_fd_sc_hd__sdfbbn_1 c331 (.CLK_N(clknet_4_2_0_clk),
    .D(net176),
    .RESET_B(net320),
    .SCD(net314),
    .SCE(net317),
    .SET_B(net306),
    .Q(net321));
 sky130_fd_sc_hd__and3_1 c332 (.A(net311),
    .B(net773),
    .C(net320),
    .X(net322));
 sky130_fd_sc_hd__and3_1 c333 (.A(net797),
    .B(net322),
    .C(net773),
    .X(net323));
 sky130_fd_sc_hd__sdfbbp_1 c334 (.CLK(clknet_4_3_0_clk),
    .D(net779),
    .RESET_B(net323),
    .SCD(net320),
    .SCE(net306),
    .SET_B(net322),
    .Q(net324));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(net324),
    .A1(net321),
    .A2(net323),
    .A3(net320),
    .S0(net305),
    .S1(net306),
    .X(net325));
 sky130_fd_sc_hd__and2_1 c336 (.A(net203),
    .B(net709),
    .X(net326));
 sky130_fd_sc_hd__and2_2 c337 (.A(net326),
    .B(net67),
    .X(net327));
 sky130_fd_sc_hd__and2_0 c338 (.A(net327),
    .B(net326),
    .X(net328));
 sky130_fd_sc_hd__and2_0 c339 (.A(net326),
    .B(net206),
    .X(net329));
 sky130_fd_sc_hd__and3_1 c34 (.A(net4),
    .B(net732),
    .C(net734),
    .X(net9));
 sky130_fd_sc_hd__and2_1 c340 (.A(net329),
    .B(net327),
    .X(net330));
 sky130_fd_sc_hd__and2_1 c341 (.A(net328),
    .B(net206),
    .X(net331));
 sky130_fd_sc_hd__and2_1 c342 (.A(net329),
    .B(net327),
    .X(net332));
 sky130_fd_sc_hd__and2_1 c343 (.A(net331),
    .B(net327),
    .X(net333));
 sky130_fd_sc_hd__sdlclkp_1 c344 (.CLK(clknet_4_9_0_clk),
    .GATE(net330),
    .SCE(net333),
    .GCLK(net334));
 sky130_fd_sc_hd__sdlclkp_2 c345 (.CLK(clknet_4_9_0_clk),
    .GATE(net326),
    .SCE(net333),
    .GCLK(net335));
 sky130_fd_sc_hd__and2_0 c346 (.A(clknet_1_1__leaf_net335),
    .B(net332),
    .X(net336));
 sky130_fd_sc_hd__and2_0 c347 (.A(net328),
    .B(clknet_1_0__leaf_net336),
    .X(net337));
 sky130_fd_sc_hd__and2_0 c348 (.A(net331),
    .B(clknet_1_0__leaf_net336),
    .X(net338));
 sky130_fd_sc_hd__and3_2 c349 (.A(net332),
    .B(net331),
    .C(net326),
    .X(net339));
 sky130_fd_sc_hd__or4bb_1 c35 (.A(net5),
    .B(net8),
    .C_N(net7),
    .D_N(net730),
    .X(net10));
 sky130_fd_sc_hd__sdfxtp_1 c350 (.CLK(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net338),
    .SCD(net339),
    .SCE(net326),
    .Q(net340));
 sky130_fd_sc_hd__dfbbn_1 c351 (.CLK_N(clknet_4_8_0_clk),
    .D(net330),
    .RESET_B(clknet_1_1__leaf_net337),
    .SET_B(clknet_1_0__leaf_net335),
    .Q(net342),
    .Q_N(net341));
 sky130_fd_sc_hd__sdfrbp_1 c352 (.CLK(clknet_4_9_0_clk),
    .D(net333),
    .RESET_B(net330),
    .SCD(clknet_1_0__leaf_net337),
    .SCE(net327),
    .Q(net344),
    .Q_N(net343));
 sky130_fd_sc_hd__dfbbn_1 c353 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net334),
    .RESET_B(net340),
    .SET_B(clknet_1_1__leaf_net338),
    .Q(net346),
    .Q_N(net345));
 sky130_fd_sc_hd__and2_0 c354 (.A(net344),
    .B(clknet_1_1__leaf_net336),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net340),
    .A1(clknet_1_0__leaf_net347),
    .A2(net341),
    .A3(clknet_1_1__leaf_net334),
    .S0(net327),
    .S1(net332),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(net345),
    .A1(net339),
    .A2(net343),
    .A3(net331),
    .S0(net709),
    .S1(net782),
    .X(net349));
 sky130_fd_sc_hd__and2_0 c357 (.A(net236),
    .B(net327),
    .X(net350));
 sky130_fd_sc_hd__and2_1 c358 (.A(net219),
    .B(net753),
    .X(net351));
 sky130_fd_sc_hd__and2_1 c359 (.A(net238),
    .B(net351),
    .X(net352));
 sky130_fd_sc_hd__and2_0 c36 (.A(net9),
    .B(net10),
    .X(net11));
 sky130_fd_sc_hd__and2_1 c360 (.A(net350),
    .B(net351),
    .X(net353));
 sky130_fd_sc_hd__sdlclkp_4 c361 (.CLK(clknet_4_10_0_clk),
    .GATE(clknet_1_1__leaf_net347),
    .SCE(net353),
    .GCLK(net354));
 sky130_fd_sc_hd__and2_2 c362 (.A(net353),
    .B(net351),
    .X(net355));
 sky130_fd_sc_hd__dfrbp_1 c363 (.CLK(clknet_4_10_0_clk),
    .D(net354),
    .RESET_B(net355),
    .Q(net357),
    .Q_N(net356));
 sky130_fd_sc_hd__and2_1 c364 (.A(net764),
    .B(net353),
    .X(net358));
 sky130_fd_sc_hd__and2_1 c365 (.A(net342),
    .B(net351),
    .X(net359));
 sky130_fd_sc_hd__dfrbp_1 c366 (.CLK(clknet_4_10_0_clk),
    .D(net352),
    .RESET_B(net355),
    .Q(net360));
 sky130_fd_sc_hd__dfrtn_1 c367 (.CLK_N(clknet_4_11_0_clk),
    .D(net339),
    .RESET_B(net358),
    .Q(net361));
 sky130_fd_sc_hd__dfrtp_1 c368 (.CLK(clknet_4_10_0_clk),
    .D(net232),
    .RESET_B(net358),
    .Q(net362));
 sky130_fd_sc_hd__or4bb_1 c369 (.A(net361),
    .B(net359),
    .C_N(net356),
    .D_N(net217),
    .X(net363));
 sky130_fd_sc_hd__a2111o_1 c37 (.A1(net11),
    .A2(net6),
    .B1(net725),
    .C1(net7),
    .D1(net730),
    .X(net12));
 sky130_fd_sc_hd__and2_0 c370 (.A(net360),
    .B(net359),
    .X(net364));
 sky130_fd_sc_hd__dfrtp_1 c371 (.CLK(clknet_4_10_0_clk),
    .D(net363),
    .RESET_B(net355),
    .Q(net365));
 sky130_fd_sc_hd__and2_1 c372 (.A(net359),
    .B(net357),
    .X(net366));
 sky130_fd_sc_hd__and2_0 c373 (.A(net364),
    .B(net365),
    .X(net367));
 sky130_fd_sc_hd__sdfbbn_1 c374 (.CLK_N(clknet_4_11_0_clk),
    .D(net366),
    .RESET_B(net355),
    .SCD(net358),
    .SCE(net339),
    .SET_B(net362),
    .Q(net369),
    .Q_N(net368));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net367),
    .A1(net353),
    .A2(net369),
    .A3(net359),
    .S0(net366),
    .S1(net355),
    .X(net370));
 sky130_fd_sc_hd__and2_0 c376 (.A(net369),
    .B(net713),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net796),
    .A1(net371),
    .A2(net366),
    .A3(net368),
    .S0(net353),
    .S1(net352),
    .X(net372));
 sky130_fd_sc_hd__buf_1 c378 (.A(net248),
    .X(net373));
 sky130_fd_sc_hd__and2_0 c379 (.A(net373),
    .B(net250),
    .X(net374));
 sky130_fd_sc_hd__and3_1 c38 (.A(net12),
    .B(net11),
    .C(net718),
    .X(net13));
 sky130_fd_sc_hd__and2_0 c380 (.A(net373),
    .B(net374),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 c381 (.A(net373),
    .X(net376));
 sky130_fd_sc_hd__and2_1 c382 (.A(net376),
    .B(net373),
    .X(net377));
 sky130_fd_sc_hd__and2_0 c383 (.A(net377),
    .B(net373),
    .X(net378));
 sky130_fd_sc_hd__and2_1 c384 (.A(net259),
    .B(net377),
    .X(net379));
 sky130_fd_sc_hd__and2_0 c385 (.A(net377),
    .B(net379),
    .X(net380));
 sky130_fd_sc_hd__and3_1 c386 (.A(net374),
    .B(net377),
    .C(net373),
    .X(net381));
 sky130_fd_sc_hd__and2_0 c387 (.A(net375),
    .B(net381),
    .X(net382));
 sky130_fd_sc_hd__and2_0 c388 (.A(net380),
    .B(net379),
    .X(net383));
 sky130_fd_sc_hd__and2_0 c389 (.A(net378),
    .B(net374),
    .X(net384));
 sky130_fd_sc_hd__or4bb_1 c39 (.A(net0),
    .B(net12),
    .C_N(net730),
    .D_N(net5),
    .X(net14));
 sky130_fd_sc_hd__and3_1 c390 (.A(net250),
    .B(net383),
    .C(net379),
    .X(net385));
 sky130_fd_sc_hd__and2_0 c391 (.A(net384),
    .B(net385),
    .X(net386));
 sky130_fd_sc_hd__and3_1 c392 (.A(net381),
    .B(net380),
    .C(net378),
    .X(net387));
 sky130_fd_sc_hd__and3_1 c393 (.A(net387),
    .B(net378),
    .C(net375),
    .X(net388));
 sky130_fd_sc_hd__and3_1 c394 (.A(net379),
    .B(net382),
    .C(net388),
    .X(net389));
 sky130_fd_sc_hd__and2_0 c395 (.A(net383),
    .B(net386),
    .X(net390));
 sky130_fd_sc_hd__dfrtp_1 c396 (.CLK(clknet_4_4_0_clk),
    .D(net376),
    .RESET_B(net390),
    .Q(net391));
 sky130_fd_sc_hd__and3_1 c397 (.A(net386),
    .B(net765),
    .C(net373),
    .X(net392));
 sky130_fd_sc_hd__dfbbp_1 c398 (.CLK(clknet_4_5_0_clk),
    .D(net392),
    .RESET_B(net390),
    .SET_B(net765),
    .Q(net394),
    .Q_N(net393));
 sky130_fd_sc_hd__buf_6 c399 (.A(net708),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c40 (.A0(net729),
    .A1(net14),
    .A2(net9),
    .A3(net7),
    .S0(net730),
    .S1(net732),
    .X(net15));
 sky130_fd_sc_hd__and2_1 c400 (.A(net385),
    .B(net395),
    .X(net396));
 sky130_fd_sc_hd__buf_1 c401 (.A(net799),
    .X(net397));
 sky130_fd_sc_hd__and2_1 c402 (.A(net395),
    .B(net388),
    .X(net398));
 sky130_fd_sc_hd__buf_1 c403 (.A(net398),
    .X(net399));
 sky130_fd_sc_hd__dfsbp_1 c404 (.CLK(clknet_4_4_0_clk),
    .D(net397),
    .SET_B(net399),
    .Q(net401),
    .Q_N(net400));
 sky130_fd_sc_hd__and2_0 c405 (.A(net395),
    .B(net397),
    .X(net402));
 sky130_fd_sc_hd__dfsbp_1 c406 (.CLK(clknet_4_5_0_clk),
    .D(net399),
    .SET_B(net397),
    .Q(net403));
 sky130_fd_sc_hd__sdfxbp_1 c407 (.CLK(clknet_4_7_0_clk),
    .D(net399),
    .SCD(net784),
    .SCE(net396),
    .Q(net405),
    .Q_N(net404));
 sky130_fd_sc_hd__and2_0 c408 (.A(net402),
    .B(net404),
    .X(net406));
 sky130_fd_sc_hd__and2_0 c409 (.A(net397),
    .B(net406),
    .X(net407));
 sky130_fd_sc_hd__and3_1 c41 (.A(net6),
    .B(net15),
    .C(net7),
    .X(net16));
 sky130_fd_sc_hd__and2_4 c410 (.A(net395),
    .B(net403),
    .X(net408));
 sky130_fd_sc_hd__and2_4 c411 (.A(net408),
    .B(net405),
    .X(net409));
 sky130_fd_sc_hd__dfstp_1 c412 (.CLK(clknet_4_4_0_clk),
    .D(net407),
    .SET_B(net399),
    .Q(net410));
 sky130_fd_sc_hd__and2_4 c413 (.A(net409),
    .B(net410),
    .X(net411));
 sky130_fd_sc_hd__and3_1 c414 (.A(net411),
    .B(net405),
    .C(net409),
    .X(net412));
 sky130_fd_sc_hd__and3_1 c415 (.A(net396),
    .B(net405),
    .C(net410),
    .X(net413));
 sky130_fd_sc_hd__sdfxbp_1 c416 (.CLK(clknet_4_6_0_clk),
    .D(net406),
    .SCD(net413),
    .SCE(net801),
    .Q(net415),
    .Q_N(net414));
 sky130_fd_sc_hd__and3_1 c417 (.A(net411),
    .B(net410),
    .C(net398),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net804),
    .A1(net416),
    .A2(net412),
    .A3(net404),
    .S0(net413),
    .S1(net411),
    .X(net417));
 sky130_fd_sc_hd__and3_1 c419 (.A(net398),
    .B(net414),
    .C(net802),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 c42 (.A(net13),
    .X(net17));
 sky130_fd_sc_hd__dfstp_1 c420 (.CLK(clknet_4_6_0_clk),
    .D(net416),
    .SET_B(net286),
    .Q(net419));
 sky130_fd_sc_hd__dfstp_1 c421 (.CLK(clknet_4_3_0_clk),
    .D(net286),
    .SET_B(net766),
    .Q(net420));
 sky130_fd_sc_hd__and2_0 c422 (.A(net419),
    .B(net272),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 c423 (.A(net420),
    .X(net422));
 sky130_fd_sc_hd__and2_0 c424 (.A(net303),
    .B(net420),
    .X(net423));
 sky130_fd_sc_hd__dfxbp_1 c425 (.CLK(clknet_4_6_0_clk),
    .D(net418),
    .Q(net425),
    .Q_N(net424));
 sky130_fd_sc_hd__and2_0 c426 (.A(net425),
    .B(net422),
    .X(net426));
 sky130_fd_sc_hd__and2_4 c427 (.A(net412),
    .B(net425),
    .X(net427));
 sky130_fd_sc_hd__and2_0 c428 (.A(net421),
    .B(net794),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 c429 (.A(net425),
    .X(net429));
 sky130_fd_sc_hd__and2_0 c43 (.A(net17),
    .B(net7),
    .X(net18));
 sky130_fd_sc_hd__and2_4 c430 (.A(net427),
    .B(net426),
    .X(net430));
 sky130_fd_sc_hd__and2_0 c431 (.A(net429),
    .B(net424),
    .X(net431));
 sky130_fd_sc_hd__dlrbn_1 c432 (.D(net430),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net428),
    .Q(net433),
    .Q_N(net432));
 sky130_fd_sc_hd__and3_1 c433 (.A(net430),
    .B(net426),
    .C(net433),
    .X(net434));
 sky130_fd_sc_hd__and2_0 c434 (.A(net401),
    .B(net429),
    .X(net435));
 sky130_fd_sc_hd__or4bb_1 c435 (.A(net427),
    .B(net435),
    .C_N(net434),
    .D_N(net432),
    .X(net436));
 sky130_fd_sc_hd__and3_1 c436 (.A(net434),
    .B(net435),
    .C(net433),
    .X(net437));
 sky130_fd_sc_hd__a2111o_1 c437 (.A1(net431),
    .A2(net436),
    .B1(net806),
    .C1(net437),
    .D1(net424),
    .X(net438));
 sky130_fd_sc_hd__or4bb_1 c438 (.A(net423),
    .B(net438),
    .C_N(net421),
    .D_N(net810),
    .X(net439));
 sky130_fd_sc_hd__sdfbbn_1 c439 (.CLK_N(clknet_4_6_0_clk),
    .D(net438),
    .RESET_B(net439),
    .SCD(net431),
    .SCE(net437),
    .SET_B(net769),
    .Q(net441),
    .Q_N(net440));
 sky130_fd_sc_hd__buf_1 c44 (.A(net14),
    .X(net19));
 sky130_fd_sc_hd__and3_1 c440 (.A(net437),
    .B(net441),
    .C(net422),
    .X(net442));
 sky130_fd_sc_hd__dfxbp_1 c441 (.CLK(clknet_4_3_0_clk),
    .D(net428),
    .Q(net444),
    .Q_N(net443));
 sky130_fd_sc_hd__buf_1 c442 (.A(net443),
    .X(net445));
 sky130_fd_sc_hd__buf_1 c443 (.A(net444),
    .X(net446));
 sky130_fd_sc_hd__and2_1 c444 (.A(net444),
    .B(net446),
    .X(net447));
 sky130_fd_sc_hd__or4bb_1 c445 (.A(net442),
    .B(net445),
    .C_N(net446),
    .D_N(net447),
    .X(net448));
 sky130_fd_sc_hd__and2_0 c446 (.A(net446),
    .B(net447),
    .X(net449));
 sky130_fd_sc_hd__and2_1 c447 (.A(net445),
    .B(net447),
    .X(net450));
 sky130_fd_sc_hd__and3_1 c448 (.A(net312),
    .B(net448),
    .C(net443),
    .X(net451));
 sky130_fd_sc_hd__or4bb_1 c449 (.A(net450),
    .B(net447),
    .C_N(net451),
    .D_N(net440),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 c45 (.A(net19),
    .X(net20));
 sky130_fd_sc_hd__and3_1 c450 (.A(net451),
    .B(net448),
    .C(net450),
    .X(net453));
 sky130_fd_sc_hd__and3_1 c451 (.A(net451),
    .B(net445),
    .C(net453),
    .X(net454));
 sky130_fd_sc_hd__and2_1 c452 (.A(net454),
    .B(net450),
    .X(net455));
 sky130_fd_sc_hd__and3_1 c453 (.A(net441),
    .B(net452),
    .C(net453),
    .X(net456));
 sky130_fd_sc_hd__and3_1 c454 (.A(net456),
    .B(net453),
    .C(net455),
    .X(net457));
 sky130_fd_sc_hd__and3_1 c455 (.A(net453),
    .B(net455),
    .C(net447),
    .X(net458));
 sky130_fd_sc_hd__and2_0 c456 (.A(net449),
    .B(net455),
    .X(net459));
 sky130_fd_sc_hd__and3_1 c457 (.A(net445),
    .B(net459),
    .C(net454),
    .X(net460));
 sky130_fd_sc_hd__or4bb_1 c458 (.A(net310),
    .B(net457),
    .C_N(net447),
    .D_N(net454),
    .X(net461));
 sky130_fd_sc_hd__and3_1 c459 (.A(net460),
    .B(net461),
    .C(net454),
    .X(net462));
 sky130_fd_sc_hd__and2_1 c46 (.A(net18),
    .B(net20),
    .X(net21));
 sky130_fd_sc_hd__and3_1 c460 (.A(net458),
    .B(net462),
    .C(net455),
    .X(net463));
 sky130_fd_sc_hd__a2111o_1 c461 (.A1(net454),
    .A2(net463),
    .B1(net451),
    .C1(net446),
    .D1(net461),
    .X(net464));
 sky130_fd_sc_hd__and2_1 c462 (.A(net464),
    .B(net793),
    .X(net465));
 sky130_fd_sc_hd__dfxtp_1 c463 (.CLK(clknet_4_12_0_clk),
    .D(net465),
    .Q(net466));
 sky130_fd_sc_hd__and2_1 c464 (.A(net448),
    .B(net781),
    .X(net467));
 sky130_fd_sc_hd__dlrbn_1 c465 (.D(net781),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net465),
    .Q(net468));
 sky130_fd_sc_hd__and2_2 c466 (.A(net327),
    .B(net711),
    .X(net469));
 sky130_fd_sc_hd__and2_1 c467 (.A(net467),
    .B(net469),
    .X(net470));
 sky130_fd_sc_hd__and2_2 c468 (.A(net450),
    .B(net469),
    .X(net744));
 sky130_fd_sc_hd__and2_1 c469 (.A(net783),
    .B(net467),
    .X(net471));
 sky130_fd_sc_hd__and3_1 c47 (.A(net21),
    .B(net18),
    .C(net20),
    .X(net22));
 sky130_fd_sc_hd__and3_1 c470 (.A(net469),
    .B(net471),
    .C(net470),
    .X(net472));
 sky130_fd_sc_hd__sdfxtp_1 c471 (.CLK(clknet_4_12_0_clk),
    .D(net465),
    .SCD(net470),
    .SCE(net744),
    .Q(net473));
 sky130_fd_sc_hd__and2_2 c472 (.A(net346),
    .B(net744),
    .X(net474));
 sky130_fd_sc_hd__sdfxtp_1 c473 (.CLK(clknet_4_11_0_clk),
    .D(net470),
    .SCD(net474),
    .SCE(net472),
    .Q(net475));
 sky130_fd_sc_hd__sdfxtp_1 c474 (.CLK(clknet_4_14_0_clk),
    .D(net781),
    .SCD(net776),
    .SCE(net474),
    .Q(net476));
 sky130_fd_sc_hd__sdfrbp_1 c475 (.CLK(clknet_4_14_0_clk),
    .D(net761),
    .RESET_B(net474),
    .SCD(net339),
    .SCE(net469),
    .Q(net477));
 sky130_fd_sc_hd__sdfrtn_1 c476 (.CLK_N(clknet_4_9_0_clk),
    .D(net447),
    .RESET_B(net760),
    .SCD(net469),
    .SCE(net474),
    .Q(net478));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net478),
    .A1(net469),
    .A2(net476),
    .A3(net466),
    .S0(net744),
    .S1(net712),
    .X(net479));
 sky130_fd_sc_hd__dfbbn_1 c478 (.CLK_N(clknet_4_14_0_clk),
    .D(net479),
    .RESET_B(net471),
    .SET_B(net467),
    .Q(net481),
    .Q_N(net480));
 sky130_fd_sc_hd__sdfrtp_1 c479 (.CLK(clknet_4_14_0_clk),
    .D(net471),
    .RESET_B(net761),
    .SCD(net481),
    .SCE(net479),
    .Q(net482));
 sky130_fd_sc_hd__and2_0 c48 (.A(net13),
    .B(net22),
    .X(net23));
 sky130_fd_sc_hd__sdfrtp_1 c480 (.CLK(clknet_4_11_0_clk),
    .D(net777),
    .RESET_B(net471),
    .SCD(net478),
    .SCE(net479),
    .Q(net483));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net798),
    .A1(net809),
    .A2(net480),
    .A3(net478),
    .S0(net339),
    .S1(net469),
    .X(net484));
 sky130_fd_sc_hd__sdfbbp_1 c482 (.CLK(clknet_4_14_0_clk),
    .D(net481),
    .RESET_B(net479),
    .SCD(net761),
    .SCE(net474),
    .SET_B(net762),
    .Q(net742),
    .Q_N(net485));
 sky130_fd_sc_hd__dlrbp_1 c487 (.D(net472),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net485),
    .Q(net752),
    .Q_N(net486));
 sky130_fd_sc_hd__dlrbp_1 c488 (.D(net372),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net744),
    .Q(net488),
    .Q_N(net487));
 sky130_fd_sc_hd__and2_0 c489 (.A(net214),
    .B(net487),
    .X(net489));
 sky130_fd_sc_hd__and2_0 c49 (.A(net20),
    .B(net17),
    .X(net24));
 sky130_fd_sc_hd__dlrtn_1 c490 (.D(net489),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net372),
    .Q(net490));
 sky130_fd_sc_hd__and2_0 c491 (.A(net752),
    .B(net490),
    .X(net491));
 sky130_fd_sc_hd__and2_0 c492 (.A(net490),
    .B(net491),
    .X(net492));
 sky130_fd_sc_hd__and2_0 c493 (.A(net488),
    .B(net486),
    .X(net493));
 sky130_fd_sc_hd__and2_1 c494 (.A(net490),
    .B(net492),
    .X(net494));
 sky130_fd_sc_hd__and2_0 c495 (.A(net491),
    .B(net494),
    .X(net749));
 sky130_fd_sc_hd__and3_1 c496 (.A(net488),
    .B(net494),
    .C(net485),
    .X(net748));
 sky130_fd_sc_hd__and2_0 c497 (.A(net749),
    .B(net494),
    .X(net741));
 sky130_fd_sc_hd__and2_0 c498 (.A(net491),
    .B(net748),
    .X(net750));
 sky130_fd_sc_hd__and3_1 c499 (.A(net492),
    .B(net489),
    .C(net750),
    .X(net747));
 sky130_fd_sc_hd__and3_1 c50 (.A(net7),
    .B(net23),
    .C(net20),
    .X(net25));
 sky130_fd_sc_hd__and3_1 c500 (.A(net493),
    .B(net748),
    .C(net747),
    .X(net745));
 sky130_fd_sc_hd__and3_1 c501 (.A(net489),
    .B(net492),
    .C(net750),
    .X(net740));
 sky130_fd_sc_hd__and3_1 c502 (.A(net494),
    .B(net745),
    .C(net747),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c503 (.A(net493),
    .B(net495),
    .C(net740),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 c504 (.A(net389),
    .X(net496));
 sky130_fd_sc_hd__dfxtp_1 c505 (.CLK(clknet_4_5_0_clk),
    .D(net496),
    .Q(net497));
 sky130_fd_sc_hd__clkbuf_1 c506 (.A(net497),
    .X(net498));
 sky130_fd_sc_hd__and2_2 c507 (.A(net498),
    .B(net385),
    .X(net499));
 sky130_fd_sc_hd__and2_0 c508 (.A(net498),
    .B(net497),
    .X(net500));
 sky130_fd_sc_hd__and2_1 c509 (.A(net498),
    .B(net785),
    .X(net501));
 sky130_fd_sc_hd__and2_0 c51 (.A(net19),
    .B(net20),
    .X(net26));
 sky130_fd_sc_hd__and3_1 c510 (.A(net497),
    .B(net501),
    .C(net499),
    .X(net502));
 sky130_fd_sc_hd__and2_0 c511 (.A(net501),
    .B(net500),
    .X(net503));
 sky130_fd_sc_hd__dlrtn_1 c512 (.D(net502),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net786),
    .Q(net504));
 sky130_fd_sc_hd__and3_1 c513 (.A(net503),
    .B(net499),
    .C(net500),
    .X(net505));
 sky130_fd_sc_hd__dlrtn_1 c514 (.D(net504),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net505),
    .Q(net506));
 sky130_fd_sc_hd__dlrtp_1 c515 (.D(net500),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net502),
    .Q(net507));
 sky130_fd_sc_hd__dfbbn_1 c516 (.CLK_N(clknet_4_5_0_clk),
    .D(net770),
    .RESET_B(net771),
    .SET_B(net502),
    .Q(net509),
    .Q_N(net508));
 sky130_fd_sc_hd__and2_1 c517 (.A(net389),
    .B(net767),
    .X(net510));
 sky130_fd_sc_hd__dfbbp_1 c518 (.CLK(clknet_4_5_0_clk),
    .D(net509),
    .RESET_B(net510),
    .SET_B(net767),
    .Q(net512),
    .Q_N(net511));
 sky130_fd_sc_hd__or4bb_1 c519 (.A(net512),
    .B(net499),
    .C_N(net508),
    .D_N(net507),
    .X(net513));
 sky130_fd_sc_hd__and2_1 c52 (.A(net24),
    .B(net19),
    .X(net27));
 sky130_fd_sc_hd__sdfxbp_1 c520 (.CLK(clknet_4_5_0_clk),
    .D(net388),
    .SCD(net513),
    .SCE(net512),
    .Q(net514));
 sky130_fd_sc_hd__sdfxbp_1 c521 (.CLK(clknet_4_5_0_clk),
    .D(net774),
    .SCD(net513),
    .SCE(net767),
    .Q(net515));
 sky130_fd_sc_hd__sdfxtp_1 c522 (.CLK(clknet_4_5_0_clk),
    .D(net510),
    .SCD(net505),
    .SCE(net513),
    .Q(net516));
 sky130_fd_sc_hd__sdfrtp_1 c523 (.CLK(clknet_4_5_0_clk),
    .D(net775),
    .RESET_B(net510),
    .SCD(net505),
    .SCE(net511),
    .Q(net517));
 sky130_fd_sc_hd__and2_1 c524 (.A(net517),
    .B(net515),
    .X(net518));
 sky130_fd_sc_hd__and2_1 c525 (.A(net518),
    .B(net714),
    .X(net519));
 sky130_fd_sc_hd__dlrtp_1 c526 (.D(net519),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net416),
    .Q(net520));
 sky130_fd_sc_hd__and2_0 c527 (.A(net520),
    .B(net519),
    .X(net521));
 sky130_fd_sc_hd__and2_0 c528 (.A(net518),
    .B(net521),
    .X(net522));
 sky130_fd_sc_hd__and2_0 c529 (.A(net520),
    .B(net519),
    .X(net523));
 sky130_fd_sc_hd__and2_0 c53 (.A(net25),
    .B(net27),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c530 (.A(net275),
    .B(net520),
    .X(net524));
 sky130_fd_sc_hd__and2_0 c531 (.A(net519),
    .B(net520),
    .X(net525));
 sky130_fd_sc_hd__and2_1 c532 (.A(net521),
    .B(net523),
    .X(net526));
 sky130_fd_sc_hd__and2_0 c533 (.A(net266),
    .B(net518),
    .X(net527));
 sky130_fd_sc_hd__sdfxtp_1 c534 (.CLK(clknet_4_7_0_clk),
    .D(net524),
    .SCD(net526),
    .SCE(net805),
    .Q(net528));
 sky130_fd_sc_hd__and3_1 c535 (.A(net526),
    .B(net525),
    .C(net521),
    .X(net529));
 sky130_fd_sc_hd__and3_2 c536 (.A(net520),
    .B(net528),
    .C(net525),
    .X(net530));
 sky130_fd_sc_hd__sdfbbn_1 c537 (.CLK_N(clknet_4_7_0_clk),
    .D(net522),
    .RESET_B(net527),
    .SCD(net530),
    .SCE(net520),
    .SET_B(net418),
    .Q(net531));
 sky130_fd_sc_hd__and3_1 c538 (.A(net527),
    .B(net530),
    .C(net523),
    .X(net532));
 sky130_fd_sc_hd__and3_1 c539 (.A(net529),
    .B(net531),
    .C(net530),
    .X(net533));
 sky130_fd_sc_hd__a2111o_1 c54 (.A1(net20),
    .A2(net26),
    .B1(net28),
    .C1(net21),
    .D1(net27),
    .X(net29));
 sky130_fd_sc_hd__and3_1 c540 (.A(net532),
    .B(net529),
    .C(net520),
    .X(net534));
 sky130_fd_sc_hd__and3_1 c541 (.A(net408),
    .B(net526),
    .C(net530),
    .X(net535));
 sky130_fd_sc_hd__and3_1 c542 (.A(net525),
    .B(net528),
    .C(net535),
    .X(net536));
 sky130_fd_sc_hd__and2_0 c543 (.A(net523),
    .B(net536),
    .X(net537));
 sky130_fd_sc_hd__and2_0 c544 (.A(net537),
    .B(net535),
    .X(net538));
 sky130_fd_sc_hd__and3_1 c545 (.A(net538),
    .B(net534),
    .C(net537),
    .X(net539));
 sky130_fd_sc_hd__and2_1 c546 (.A(net437),
    .B(net499),
    .X(net540));
 sky130_fd_sc_hd__dfxtp_1 c547 (.CLK(clknet_4_12_0_clk),
    .D(net540),
    .Q(net541));
 sky130_fd_sc_hd__dlclkp_1 c548 (.CLK(clknet_4_6_0_clk),
    .GATE(net540),
    .GCLK(net542));
 sky130_fd_sc_hd__dlrtp_1 c549 (.D(net416),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(clknet_1_0__leaf_net542),
    .Q(net543));
 sky130_fd_sc_hd__and3_1 c55 (.A(net28),
    .B(net27),
    .C(net21),
    .X(net30));
 sky130_fd_sc_hd__edfxbp_1 c550 (.CLK(clknet_4_6_0_clk),
    .D(net540),
    .DE(net499),
    .Q(net544));
 sky130_fd_sc_hd__and2_0 c551 (.A(net543),
    .B(clknet_1_0__leaf_net542),
    .X(net545));
 sky130_fd_sc_hd__and3_1 c552 (.A(net544),
    .B(clknet_1_0__leaf_net545),
    .C(net518),
    .X(net546));
 sky130_fd_sc_hd__and2_0 c553 (.A(clknet_1_1__leaf_net542),
    .B(clknet_1_1__leaf_net545),
    .X(net547));
 sky130_fd_sc_hd__and3_1 c554 (.A(net442),
    .B(net543),
    .C(clknet_1_0__leaf_net542),
    .X(net548));
 sky130_fd_sc_hd__and2_0 c555 (.A(net546),
    .B(clknet_1_0__leaf_net542),
    .X(net549));
 sky130_fd_sc_hd__and3_1 c556 (.A(clknet_1_0__leaf_net547),
    .B(clknet_1_0__leaf_net548),
    .C(clknet_1_1__leaf_net542),
    .X(net550));
 sky130_fd_sc_hd__and2_0 c557 (.A(clknet_1_0__leaf_net549),
    .B(clknet_1_0__leaf_net545),
    .X(net551));
 sky130_fd_sc_hd__and2_0 c558 (.A(clknet_1_1__leaf_net551),
    .B(clknet_1_1__leaf_net547),
    .X(net552));
 sky130_fd_sc_hd__and2_4 c559 (.A(clknet_1_1__leaf_net548),
    .B(net528),
    .X(net553));
 sky130_fd_sc_hd__a2111o_1 c56 (.A1(net23),
    .A2(net30),
    .B1(net25),
    .C1(net27),
    .D1(net20),
    .X(net31));
 sky130_fd_sc_hd__and2_0 c560 (.A(clknet_1_0__leaf_net548),
    .B(clknet_1_0__leaf_net547),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c561 (.A(clknet_1_0__leaf_net554),
    .B(clknet_1_1__leaf_net549),
    .C(clknet_1_0__leaf_net551),
    .X(net555));
 sky130_fd_sc_hd__a2111o_1 c562 (.A1(net543),
    .A2(clknet_1_0__leaf_net555),
    .B1(clknet_1_0__leaf_net554),
    .C1(net530),
    .D1(clknet_1_0__leaf_net548),
    .X(net556));
 sky130_fd_sc_hd__and3_1 c563 (.A(clknet_1_1__leaf_net555),
    .B(clknet_1_0__leaf_net545),
    .C(clknet_1_0__leaf_net551),
    .X(net557));
 sky130_fd_sc_hd__and3_1 c564 (.A(clknet_1_0__leaf_net557),
    .B(clknet_1_0__leaf_net555),
    .C(clknet_1_1__leaf_net554),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net530),
    .A1(clknet_1_0__leaf_net549),
    .A2(clknet_1_0__leaf_net557),
    .A3(clknet_1_1__leaf_net542),
    .S0(clknet_1_0__leaf_net556),
    .S1(clknet_1_1__leaf_net548),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net558),
    .A1(net559),
    .A2(clknet_1_1__leaf_net553),
    .A3(clknet_1_1__leaf_net557),
    .S0(clknet_1_1__leaf_net548),
    .S1(clknet_1_1__leaf_net542),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_1 c567 (.A(net464),
    .X(net561));
 sky130_fd_sc_hd__and2_4 c568 (.A(clknet_1_0__leaf_net553),
    .B(clknet_1_1__leaf_net545),
    .X(net562));
 sky130_fd_sc_hd__buf_1 c569 (.A(net550),
    .X(net563));
 sky130_fd_sc_hd__or4bb_1 c57 (.A(net31),
    .B(net30),
    .C_N(net29),
    .D_N(net28),
    .X(net32));
 sky130_fd_sc_hd__dlclkp_2 c570 (.CLK(clknet_4_12_0_clk),
    .GATE(net561),
    .GCLK(net564));
 sky130_fd_sc_hd__and2_4 c571 (.A(net562),
    .B(clknet_1_1__leaf_net564),
    .X(net565));
 sky130_fd_sc_hd__and2_0 c572 (.A(clknet_1_0__leaf_net565),
    .B(clknet_1_1__leaf_net563),
    .X(net566));
 sky130_fd_sc_hd__and2_4 c573 (.A(clknet_1_0__leaf_net565),
    .B(net446),
    .X(net567));
 sky130_fd_sc_hd__and2_0 c574 (.A(clknet_1_0__leaf_net567),
    .B(net464),
    .X(net568));
 sky130_fd_sc_hd__edfxtp_1 c575 (.CLK(clknet_4_12_0_clk),
    .D(net568),
    .DE(clknet_1_1__leaf_net565),
    .Q(net569));
 sky130_fd_sc_hd__and2_0 c576 (.A(net569),
    .B(clknet_1_1__leaf_net565),
    .X(net754));
 sky130_fd_sc_hd__sdlclkp_1 c577 (.CLK(clknet_4_12_0_clk),
    .GATE(net561),
    .SCE(net450),
    .GCLK(net570));
 sky130_fd_sc_hd__and2_4 c578 (.A(clknet_1_0__leaf_net565),
    .B(clknet_1_0__leaf_net564),
    .X(net571));
 sky130_fd_sc_hd__and2_0 c579 (.A(clknet_1_0__leaf_net571),
    .B(clknet_1_0__leaf_net565),
    .X(net572));
 sky130_fd_sc_hd__or4bb_1 c58 (.A(net22),
    .B(net24),
    .C_N(net27),
    .D_N(net30),
    .X(net33));
 sky130_fd_sc_hd__and3_1 c580 (.A(net437),
    .B(net569),
    .C(net452),
    .X(net573));
 sky130_fd_sc_hd__and2_0 c581 (.A(net570),
    .B(clknet_1_1__leaf_net571),
    .X(net574));
 sky130_fd_sc_hd__and3_1 c582 (.A(clknet_1_1__leaf_net567),
    .B(clknet_1_0__leaf_net571),
    .C(clknet_1_0__leaf_net563),
    .X(net575));
 sky130_fd_sc_hd__and2_0 c583 (.A(net541),
    .B(clknet_1_0__leaf_net575),
    .X(net576));
 sky130_fd_sc_hd__and3_1 c584 (.A(net576),
    .B(clknet_1_0__leaf_net575),
    .C(clknet_1_0__leaf_net564),
    .X(net577));
 sky130_fd_sc_hd__or4bb_1 c585 (.A(net573),
    .B(net566),
    .C_N(clknet_1_0__leaf_net577),
    .D_N(clknet_1_0__leaf_net575),
    .X(net578));
 sky130_fd_sc_hd__and2_0 c586 (.A(net572),
    .B(net578),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net574),
    .A1(net579),
    .A2(clknet_1_0__leaf_net577),
    .A3(clknet_1_1__leaf_net575),
    .S0(clknet_1_1__leaf_net545),
    .S1(clknet_1_1__leaf_net565),
    .X(net580));
 sky130_fd_sc_hd__buf_6 c588 (.A(clknet_1_1__leaf_net575),
    .X(net581));
 sky130_fd_sc_hd__and2_0 c589 (.A(net477),
    .B(clknet_1_0__leaf_net581),
    .X(net582));
 sky130_fd_sc_hd__and3_2 c59 (.A(net32),
    .B(net31),
    .C(net30),
    .X(net34));
 sky130_fd_sc_hd__buf_6 c590 (.A(clknet_1_0__leaf_net581),
    .X(net583));
 sky130_fd_sc_hd__and2_4 c591 (.A(clknet_1_0__leaf_net583),
    .B(clknet_1_0__leaf_net581),
    .X(net584));
 sky130_fd_sc_hd__and2_0 c592 (.A(clknet_1_0__leaf_net581),
    .B(clknet_1_0__leaf_net584),
    .X(net585));
 sky130_fd_sc_hd__and2_0 c593 (.A(net585),
    .B(clknet_1_0__leaf_net584),
    .X(net586));
 sky130_fd_sc_hd__sdlclkp_2 c594 (.CLK(clknet_4_15_0_clk),
    .GATE(clknet_1_1__leaf_net556),
    .SCE(clknet_1_0__leaf_net586),
    .GCLK(net587));
 sky130_fd_sc_hd__sdfxtp_1 c595 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_0__leaf_net584),
    .SCD(clknet_1_0__leaf_net586),
    .SCE(clknet_1_0__leaf_net587),
    .Q(net588));
 sky130_fd_sc_hd__and2_4 c596 (.A(clknet_1_0__leaf_net583),
    .B(clknet_1_0__leaf_net587),
    .X(net589));
 sky130_fd_sc_hd__sdlclkp_4 c597 (.CLK(clknet_4_15_0_clk),
    .GATE(clknet_1_1__leaf_net586),
    .SCE(clknet_1_1__leaf_net589),
    .GCLK(net590));
 sky130_fd_sc_hd__and3_1 c598 (.A(net588),
    .B(clknet_1_1__leaf_net589),
    .C(clknet_1_1__leaf_net587),
    .X(net591));
 sky130_fd_sc_hd__and3_1 c599 (.A(net582),
    .B(clknet_1_0__leaf_net587),
    .C(clknet_1_0__leaf_net589),
    .X(net743));
 sky130_fd_sc_hd__or4bb_1 c60 (.A(net30),
    .B(net33),
    .C_N(net32),
    .D_N(net34),
    .X(net35));
 sky130_fd_sc_hd__and3_1 c600 (.A(clknet_1_0__leaf_net589),
    .B(clknet_1_0__leaf_net743),
    .C(clknet_1_0__leaf_net590),
    .X(net592));
 sky130_fd_sc_hd__and3_1 c601 (.A(clknet_1_1__leaf_net584),
    .B(clknet_1_0__leaf_net743),
    .C(clknet_1_1__leaf_net587),
    .X(net593));
 sky130_fd_sc_hd__and3_1 c602 (.A(clknet_1_1__leaf_net584),
    .B(clknet_1_1__leaf_net589),
    .C(clknet_1_1__leaf_net590),
    .X(net594));
 sky130_fd_sc_hd__and3_1 c603 (.A(clknet_1_0__leaf_net594),
    .B(net591),
    .C(clknet_1_0__leaf_net590),
    .X(net595));
 sky130_fd_sc_hd__dfbbn_1 c604 (.CLK_N(clknet_4_14_0_clk),
    .D(net592),
    .RESET_B(net595),
    .SET_B(clknet_1_1__leaf_net587),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__and2_0 c605 (.A(clknet_1_1__leaf_net583),
    .B(net597),
    .X(net598));
 sky130_fd_sc_hd__and3_1 c606 (.A(net598),
    .B(net597),
    .C(clknet_1_0__leaf_net594),
    .X(net599));
 sky130_fd_sc_hd__dfbbn_1 c607 (.CLK_N(clknet_4_14_0_clk),
    .D(net599),
    .RESET_B(net593),
    .SET_B(net596),
    .Q(net600));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(clknet_1_1__leaf_net581),
    .A1(net600),
    .A2(clknet_1_1__leaf_net594),
    .A3(clknet_1_1__leaf_net577),
    .S0(clknet_1_1__leaf_net590),
    .S1(clknet_1_1__leaf_net587),
    .X(net751));
 sky130_fd_sc_hd__or4bb_1 c61 (.A(net27),
    .B(net35),
    .C_N(net34),
    .D_N(net30),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net36),
    .A1(net29),
    .A2(net35),
    .A3(net30),
    .S0(net34),
    .S1(net20),
    .X(net37));
 sky130_fd_sc_hd__dfrbp_1 c63 (.CLK(clknet_4_0_0_clk),
    .D(net34),
    .RESET_B(net37),
    .Q(net39),
    .Q_N(net38));
 sky130_fd_sc_hd__buf_1 c630 (.A(net518),
    .X(net601));
 sky130_fd_sc_hd__buf_1 c631 (.A(net601),
    .X(net602));
 sky130_fd_sc_hd__and2_0 c632 (.A(net601),
    .B(net602),
    .X(net603));
 sky130_fd_sc_hd__buf_1 c633 (.A(net602),
    .X(net604));
 sky130_fd_sc_hd__and2_1 c634 (.A(net604),
    .B(net601),
    .X(net605));
 sky130_fd_sc_hd__and2_1 c635 (.A(net603),
    .B(net605),
    .X(net606));
 sky130_fd_sc_hd__and2_0 c636 (.A(net605),
    .B(net602),
    .X(net607));
 sky130_fd_sc_hd__and3_1 c637 (.A(net607),
    .B(net606),
    .C(net604),
    .X(net608));
 sky130_fd_sc_hd__and2_1 c638 (.A(net499),
    .B(net605),
    .X(net609));
 sky130_fd_sc_hd__dfrbp_1 c639 (.CLK(clknet_4_7_0_clk),
    .D(net609),
    .RESET_B(net606),
    .Q(net610));
 sky130_fd_sc_hd__buf_1 c64 (.A(net39),
    .X(net40));
 sky130_fd_sc_hd__and2_1 c640 (.A(net607),
    .B(net604),
    .X(net611));
 sky130_fd_sc_hd__and2_1 c641 (.A(net611),
    .B(net602),
    .X(net612));
 sky130_fd_sc_hd__and3_1 c642 (.A(net605),
    .B(net610),
    .C(net608),
    .X(net613));
 sky130_fd_sc_hd__and2_0 c643 (.A(net604),
    .B(net613),
    .X(net614));
 sky130_fd_sc_hd__and2_0 c644 (.A(net606),
    .B(net612),
    .X(net615));
 sky130_fd_sc_hd__and2_0 c645 (.A(net613),
    .B(net606),
    .X(net616));
 sky130_fd_sc_hd__sdfbbn_1 c646 (.CLK_N(clknet_4_7_0_clk),
    .D(net602),
    .RESET_B(net612),
    .SCD(net616),
    .SCE(net611),
    .SET_B(net609),
    .Q(net618),
    .Q_N(net617));
 sky130_fd_sc_hd__and2_0 c647 (.A(net618),
    .B(net615),
    .X(net619));
 sky130_fd_sc_hd__and3_1 c648 (.A(net614),
    .B(net611),
    .C(net617),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net620),
    .A1(net616),
    .A2(net611),
    .A3(net608),
    .S0(net601),
    .S1(net613),
    .X(net621));
 sky130_fd_sc_hd__dfrbp_1 c65 (.CLK(clknet_4_0_0_clk),
    .D(net40),
    .RESET_B(net37),
    .Q(net42),
    .Q_N(net41));
 sky130_fd_sc_hd__and3_1 c650 (.A(net621),
    .B(net620),
    .C(net611),
    .X(net622));
 sky130_fd_sc_hd__and2_1 c651 (.A(net622),
    .B(net608),
    .X(net623));
 sky130_fd_sc_hd__and2_0 c652 (.A(net623),
    .B(net530),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 c653 (.A(net612),
    .X(net625));
 sky130_fd_sc_hd__and2_0 c654 (.A(net625),
    .B(net624),
    .X(net626));
 sky130_fd_sc_hd__and2_1 c655 (.A(net624),
    .B(net623),
    .X(net627));
 sky130_fd_sc_hd__and2_0 c656 (.A(net625),
    .B(net612),
    .X(net628));
 sky130_fd_sc_hd__and2_1 c657 (.A(net626),
    .B(net623),
    .X(net629));
 sky130_fd_sc_hd__and2_0 c658 (.A(net619),
    .B(net624),
    .X(net630));
 sky130_fd_sc_hd__and2_0 c659 (.A(net630),
    .B(net627),
    .X(net631));
 sky130_fd_sc_hd__and2_1 c66 (.A(net41),
    .B(net40),
    .X(net43));
 sky130_fd_sc_hd__and2_0 c660 (.A(net631),
    .B(net625),
    .X(net632));
 sky130_fd_sc_hd__and3_1 c661 (.A(net533),
    .B(net630),
    .C(net631),
    .X(net633));
 sky130_fd_sc_hd__and3_1 c662 (.A(net629),
    .B(net631),
    .C(net633),
    .X(net634));
 sky130_fd_sc_hd__and3_1 c663 (.A(net627),
    .B(net634),
    .C(net633),
    .X(net635));
 sky130_fd_sc_hd__and3_1 c664 (.A(net539),
    .B(net634),
    .C(net635),
    .X(net636));
 sky130_fd_sc_hd__dfbbp_1 c665 (.CLK(clknet_4_7_0_clk),
    .D(net636),
    .RESET_B(net635),
    .SET_B(net633),
    .Q(net637));
 sky130_fd_sc_hd__a2111o_1 c666 (.A1(net628),
    .A2(net635),
    .B1(net623),
    .C1(net627),
    .D1(net633),
    .X(net638));
 sky130_fd_sc_hd__or4bb_1 c667 (.A(net608),
    .B(net637),
    .C_N(net638),
    .D_N(net635),
    .X(net639));
 sky130_fd_sc_hd__and2_0 c668 (.A(net632),
    .B(net638),
    .X(net640));
 sky130_fd_sc_hd__sdfbbp_1 c669 (.CLK(clknet_4_13_0_clk),
    .D(net640),
    .RESET_B(net633),
    .SCD(net638),
    .SCE(net627),
    .SET_B(net625),
    .Q(net641));
 sky130_fd_sc_hd__and2_2 c67 (.A(net40),
    .B(net43),
    .X(net44));
 sky130_fd_sc_hd__sdfsbp_1 c670 (.CLK(clknet_4_13_0_clk),
    .D(net633),
    .SCD(net639),
    .SCE(net632),
    .SET_B(net629),
    .Q(net642));
 sky130_fd_sc_hd__and3_1 c671 (.A(net807),
    .B(net768),
    .C(net638),
    .X(net643));
 sky130_fd_sc_hd__dlclkp_4 c672 (.CLK(clknet_4_13_0_clk),
    .GATE(net643),
    .GCLK(net644));
 sky130_fd_sc_hd__and2_0 c673 (.A(net560),
    .B(net625),
    .X(net645));
 sky130_fd_sc_hd__dlxbn_1 c674 (.D(net643),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net646));
 sky130_fd_sc_hd__buf_1 c675 (.A(net625),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 c676 (.A(net647),
    .X(net648));
 sky130_fd_sc_hd__and3_1 c677 (.A(net645),
    .B(net648),
    .C(net625),
    .X(net649));
 sky130_fd_sc_hd__and2_0 c678 (.A(clknet_1_0__leaf_net545),
    .B(net622),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 c679 (.A(net648),
    .X(net651));
 sky130_fd_sc_hd__dfrtn_1 c68 (.CLK_N(clknet_4_0_0_clk),
    .D(net37),
    .RESET_B(net43),
    .Q(net45));
 sky130_fd_sc_hd__and2_0 c680 (.A(net648),
    .B(clknet_1_0__leaf_net649),
    .X(net652));
 sky130_fd_sc_hd__and2_0 c681 (.A(net552),
    .B(clknet_1_0__leaf_net644),
    .X(net653));
 sky130_fd_sc_hd__sdfxbp_1 c682 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_0__leaf_net649),
    .SCD(net643),
    .SCE(net648),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__and2_0 c683 (.A(clknet_1_1__leaf_net644),
    .B(clknet_1_1__leaf_net649),
    .X(net656));
 sky130_fd_sc_hd__or4bb_1 c684 (.A(net650),
    .B(clknet_1_0__leaf_net653),
    .C_N(clknet_1_0__leaf_net644),
    .D_N(net654),
    .X(net657));
 sky130_fd_sc_hd__and3_1 c685 (.A(net646),
    .B(clknet_1_1__leaf_net653),
    .C(clknet_1_0__leaf_net656),
    .X(net658));
 sky130_fd_sc_hd__a2111o_1 c686 (.A1(net652),
    .A2(net647),
    .B1(net648),
    .C1(clknet_1_0__leaf_net657),
    .D1(clknet_1_1__leaf_net545),
    .X(net659));
 sky130_fd_sc_hd__and3_1 c687 (.A(clknet_1_1__leaf_net657),
    .B(net647),
    .C(net655),
    .X(net660));
 sky130_fd_sc_hd__and2_0 c688 (.A(net651),
    .B(clknet_1_0__leaf_net660),
    .X(net661));
 sky130_fd_sc_hd__or4bb_1 c689 (.A(clknet_1_1__leaf_net660),
    .B(clknet_1_0__leaf_net661),
    .C_N(clknet_1_1__leaf_net656),
    .D_N(net648),
    .X(net662));
 sky130_fd_sc_hd__and2_0 c69 (.A(net44),
    .B(net40),
    .X(net46));
 sky130_fd_sc_hd__or4bb_1 c690 (.A(clknet_1_0__leaf_net656),
    .B(net658),
    .C_N(clknet_1_1__leaf_net660),
    .D_N(clknet_1_0__leaf_net661),
    .X(net663));
 sky130_fd_sc_hd__and3_1 c691 (.A(clknet_1_1__leaf_net661),
    .B(net662),
    .C(clknet_1_1__leaf_net660),
    .X(net664));
 sky130_fd_sc_hd__sdfbbn_1 c692 (.CLK_N(clknet_4_13_0_clk),
    .D(net655),
    .RESET_B(net664),
    .SCD(net663),
    .SCE(clknet_1_0__leaf_net660),
    .SET_B(net648),
    .Q(net665));
 sky130_fd_sc_hd__dlxbn_1 c693 (.D(net580),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net666));
 sky130_fd_sc_hd__buf_1 c694 (.A(net452),
    .X(net667));
 sky130_fd_sc_hd__and2_0 c695 (.A(clknet_1_1__leaf_net577),
    .B(net667),
    .X(net668));
 sky130_fd_sc_hd__and2_1 c696 (.A(net665),
    .B(net667),
    .X(net669));
 sky130_fd_sc_hd__and2_0 c697 (.A(net669),
    .B(clknet_1_1__leaf_net575),
    .X(net670));
 sky130_fd_sc_hd__and2_0 c698 (.A(clknet_1_1__leaf_net668),
    .B(net667),
    .X(net671));
 sky130_fd_sc_hd__dfrbp_1 c699 (.CLK(clknet_4_13_0_clk),
    .D(net666),
    .RESET_B(net643),
    .Q(net673),
    .Q_N(net672));
 sky130_fd_sc_hd__dfrtp_1 c70 (.CLK(clknet_4_0_0_clk),
    .D(net43),
    .RESET_B(net37),
    .Q(net47));
 sky130_fd_sc_hd__and2_1 c700 (.A(net667),
    .B(net672),
    .X(net674));
 sky130_fd_sc_hd__and2_0 c701 (.A(net674),
    .B(net669),
    .X(net675));
 sky130_fd_sc_hd__and2_0 c702 (.A(net673),
    .B(net669),
    .X(net676));
 sky130_fd_sc_hd__and2_0 c703 (.A(clknet_1_0__leaf_net653),
    .B(net674),
    .X(net677));
 sky130_fd_sc_hd__and2_0 c704 (.A(net669),
    .B(clknet_1_0__leaf_net670),
    .X(net678));
 sky130_fd_sc_hd__and2_0 c705 (.A(clknet_1_0__leaf_net668),
    .B(clknet_1_0__leaf_net678),
    .X(net679));
 sky130_fd_sc_hd__and2_0 c706 (.A(net679),
    .B(clknet_1_0__leaf_net668),
    .X(net680));
 sky130_fd_sc_hd__dfrtn_1 c707 (.CLK_N(clknet_4_14_0_clk),
    .D(net680),
    .RESET_B(clknet_1_0__leaf_net678),
    .Q(net681));
 sky130_fd_sc_hd__and2_1 c708 (.A(net676),
    .B(net673),
    .X(net682));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net671),
    .A1(net675),
    .A2(net682),
    .A3(net674),
    .S0(net669),
    .S1(net672),
    .X(net683));
 sky130_fd_sc_hd__and3_1 c71 (.A(net42),
    .B(net47),
    .C(net46),
    .X(net48));
 sky130_fd_sc_hd__or4bb_1 c710 (.A(net681),
    .B(clknet_1_1__leaf_net678),
    .C_N(net682),
    .D_N(clknet_1_0__leaf_net670),
    .X(net684));
 sky130_fd_sc_hd__a2111o_1 c711 (.A1(net659),
    .A2(net684),
    .B1(net682),
    .C1(net530),
    .D1(net674),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net667),
    .A1(net683),
    .A2(net681),
    .A3(clknet_1_1__leaf_net668),
    .S0(net682),
    .S1(net674),
    .X(net686));
 sky130_fd_sc_hd__sdfxbp_1 c713 (.CLK(clknet_4_15_0_clk),
    .D(net682),
    .SCD(net685),
    .SCE(net788),
    .Q(net687));
 sky130_fd_sc_hd__dfrtp_1 c714 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_0__leaf_net751),
    .RESET_B(clknet_1_1__leaf_net670),
    .Q(net688));
 sky130_fd_sc_hd__and3_1 c715 (.A(net763),
    .B(net687),
    .C(clknet_1_1__leaf_net743),
    .X(net689));
 sky130_fd_sc_hd__and2_1 c716 (.A(net763),
    .B(net744),
    .X(net690));
 sky130_fd_sc_hd__sdfxtp_1 c717 (.CLK(clknet_4_15_0_clk),
    .D(net677),
    .SCD(net690),
    .SCE(clknet_1_0__leaf_net689),
    .Q(net691));
 sky130_fd_sc_hd__dfrtp_1 c718 (.CLK(clknet_4_15_0_clk),
    .D(net690),
    .RESET_B(clknet_1_0__leaf_net689),
    .Q(net692));
 sky130_fd_sc_hd__dfrtp_1 c719 (.CLK(clknet_4_15_0_clk),
    .D(net791),
    .RESET_B(net690),
    .Q(net693));
 sky130_fd_sc_hd__or4bb_2 c72 (.A(net48),
    .B(net44),
    .C_N(net45),
    .D_N(net7),
    .X(net49));
 sky130_fd_sc_hd__sdfxtp_1 c720 (.CLK(clknet_4_15_0_clk),
    .D(net763),
    .SCD(net789),
    .SCE(clknet_1_0__leaf_net751),
    .Q(net694));
 sky130_fd_sc_hd__and2_0 c721 (.A(clknet_1_1__leaf_net670),
    .B(net789),
    .X(net695));
 sky130_fd_sc_hd__and3_1 c722 (.A(net693),
    .B(net694),
    .C(net692),
    .X(net696));
 sky130_fd_sc_hd__and2_0 c723 (.A(net694),
    .B(net692),
    .X(net697));
 sky130_fd_sc_hd__dfsbp_1 c724 (.CLK(clknet_4_15_0_clk),
    .D(clknet_1_1__leaf_net689),
    .SET_B(net695),
    .Q(net698));
 sky130_fd_sc_hd__and3_1 c725 (.A(net691),
    .B(net697),
    .C(net692),
    .X(net699));
 sky130_fd_sc_hd__and3_1 c726 (.A(net697),
    .B(net694),
    .C(net692),
    .X(net700));
 sky130_fd_sc_hd__and2_0 c727 (.A(net698),
    .B(net697),
    .X(net701));
 sky130_fd_sc_hd__and3_1 c728 (.A(net696),
    .B(net699),
    .C(net692),
    .X(net702));
 sky130_fd_sc_hd__and2_0 c729 (.A(net700),
    .B(net701),
    .X(net703));
 sky130_fd_sc_hd__and2_0 c73 (.A(net40),
    .B(net49),
    .X(net50));
 sky130_fd_sc_hd__and2_0 c730 (.A(net692),
    .B(net702),
    .X(net704));
 sky130_fd_sc_hd__and3_1 c731 (.A(net704),
    .B(net703),
    .C(net702));
 sky130_fd_sc_hd__and3_1 c74 (.A(net45),
    .B(net49),
    .C(net44),
    .X(net51));
 sky130_fd_sc_hd__and2_0 c75 (.A(net51),
    .B(net48),
    .X(net52));
 sky130_fd_sc_hd__or4bb_1 c76 (.A(net43),
    .B(net49),
    .C_N(net40),
    .D_N(net51),
    .X(net53));
 sky130_fd_sc_hd__and2_0 c77 (.A(net52),
    .B(net53),
    .X(net54));
 sky130_fd_sc_hd__and2_2 c78 (.A(net53),
    .B(net54),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c79 (.A(net46),
    .B(net43),
    .C(net49),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c80 (.A0(net47),
    .A1(net56),
    .A2(net52),
    .A3(net55),
    .S0(net44),
    .S1(net38),
    .X(net57));
 sky130_fd_sc_hd__a2111o_1 c81 (.A1(net50),
    .A2(net55),
    .B1(net51),
    .C1(net49),
    .D1(net43),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net39),
    .A1(net56),
    .A2(net50),
    .A3(net55),
    .S0(net49),
    .S1(net51),
    .X(net59));
 sky130_fd_sc_hd__mux4_2 c83 (.A0(net54),
    .A1(net57),
    .A2(net58),
    .A3(net59),
    .S0(net55),
    .S1(net38),
    .X(net60));
 sky130_fd_sc_hd__buf_1 c84 (.A(net60),
    .X(net61));
 sky130_fd_sc_hd__and2_1 c85 (.A(net61),
    .B(net55),
    .X(net62));
 sky130_fd_sc_hd__and2_2 c86 (.A(net61),
    .B(net60),
    .X(net63));
 sky130_fd_sc_hd__and2_0 c87 (.A(net62),
    .B(net61),
    .X(net64));
 sky130_fd_sc_hd__and2_0 c88 (.A(net64),
    .B(net63),
    .X(net65));
 sky130_fd_sc_hd__and2_0 c89 (.A(net63),
    .B(net62),
    .X(net66));
 sky130_fd_sc_hd__and2_1 c90 (.A(net62),
    .B(net63),
    .X(net67));
 sky130_fd_sc_hd__and2_1 c91 (.A(net62),
    .B(net63),
    .X(net68));
 sky130_fd_sc_hd__and3_1 c92 (.A(net65),
    .B(net755),
    .C(net68),
    .X(net69));
 sky130_fd_sc_hd__and3_1 c93 (.A(net755),
    .B(net69),
    .C(net63),
    .X(net70));
 sky130_fd_sc_hd__and2_1 c94 (.A(net63),
    .B(net69),
    .X(net71));
 sky130_fd_sc_hd__mux4_2 c95 (.A0(net71),
    .A1(net69),
    .A2(net68),
    .A3(net62),
    .S0(net63),
    .S1(net755),
    .X(net72));
 sky130_fd_sc_hd__and3_1 c96 (.A(net68),
    .B(net69),
    .C(net72),
    .X(net73));
 sky130_fd_sc_hd__and3_1 c97 (.A(net66),
    .B(net71),
    .C(net755),
    .X(net74));
 sky130_fd_sc_hd__and3_1 c98 (.A(net74),
    .B(net71),
    .C(net72),
    .X(net75));
 sky130_fd_sc_hd__a2111o_1 c99 (.A1(net70),
    .A2(net68),
    .B1(net74),
    .C1(net66),
    .D1(net755),
    .X(net76));
 sky130_fd_sc_hd__dlxbp_1 s732 (.D(net80),
    .GATE(clknet_4_2_0_clk),
    .Q(net705));
 sky130_fd_sc_hd__dlxtn_1 s733 (.D(net81),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net706));
 sky130_fd_sc_hd__dlxtn_1 s734 (.D(net277),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net707));
 sky130_fd_sc_hd__dlxtn_2 s735 (.D(net280),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net708));
 sky130_fd_sc_hd__dlxtp_1 s736 (.D(net325),
    .GATE(clknet_4_9_0_clk),
    .Q(net709));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s737 (.D(net348),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net710));
 sky130_fd_sc_hd__dfxbp_1 s738 (.CLK(clknet_4_11_0_clk),
    .D(net349),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dfxbp_1 s739 (.CLK(clknet_4_10_0_clk),
    .D(net370),
    .Q(net713));
 sky130_fd_sc_hd__dfxtp_1 s740 (.CLK(clknet_4_6_0_clk),
    .D(net417),
    .Q(net714));
 sky130_fd_sc_hd__dfxtp_1 s741 (.CLK(clknet_4_11_0_clk),
    .D(net484),
    .Q(net715));
 sky130_fd_sc_hd__dfxtp_1 s742 (.CLK(clknet_4_15_0_clk),
    .D(net686),
    .Q(net716));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in1),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in10),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in11),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in13),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in14),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in15),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in16),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in17),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in18),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in19),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in2),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in20),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in21),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in22),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in23),
    .X(net731));
 sky130_fd_sc_hd__buf_1 input16 (.A(in24),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in3),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in4),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in5),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in6),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in7),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in8),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in9),
    .X(net739));
 sky130_fd_sc_hd__buf_2 output24 (.A(net740),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output25 (.A(net741),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output26 (.A(net742),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(clknet_1_1__leaf_net743),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output28 (.A(net744),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output29 (.A(net745),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output30 (.A(net746),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output31 (.A(net747),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output32 (.A(net748),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output33 (.A(net749),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output34 (.A(net750),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(clknet_1_1__leaf_net751),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output36 (.A(net752),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output37 (.A(net753),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net754),
    .X(out8));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net67),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net644 (.A(net644),
    .X(clknet_0_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_0__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net644 (.A(clknet_0_net644),
    .X(clknet_1_1__leaf_net644));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net660 (.A(net660),
    .X(clknet_0_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_0__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_1__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net661 (.A(net661),
    .X(clknet_0_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net661 (.A(clknet_0_net661),
    .X(clknet_1_0__leaf_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net661 (.A(clknet_0_net661),
    .X(clknet_1_1__leaf_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net653 (.A(net653),
    .X(clknet_0_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_0__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_1__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net590 (.A(net590),
    .X(clknet_0_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_0__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net590 (.A(clknet_0_net590),
    .X(clknet_1_1__leaf_net590));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net751 (.A(net751),
    .X(clknet_0_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_0__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_1__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net594 (.A(net594),
    .X(clknet_0_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_0__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net594 (.A(net756),
    .X(clknet_1_1__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net587 (.A(net587),
    .X(clknet_0_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_0__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net587 (.A(clknet_0_net587),
    .X(clknet_1_1__leaf_net587));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net743 (.A(net743),
    .X(clknet_0_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net689 (.A(net689),
    .X(clknet_0_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_0__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net689 (.A(clknet_0_net689),
    .X(clknet_1_1__leaf_net689));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net589 (.A(net589),
    .X(clknet_0_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net589 (.A(net758),
    .X(clknet_1_0__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net589 (.A(clknet_0_net589),
    .X(clknet_1_1__leaf_net589));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net564 (.A(net564),
    .X(clknet_0_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_0__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net564 (.A(clknet_0_net564),
    .X(clknet_1_1__leaf_net564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net577 (.A(net577),
    .X(clknet_0_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_0__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net577 (.A(clknet_0_net577),
    .X(clknet_1_1__leaf_net577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net668 (.A(net668),
    .X(clknet_0_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_0__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net668 (.A(clknet_0_net668),
    .X(clknet_1_1__leaf_net668));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net571 (.A(net571),
    .X(clknet_0_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_0__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net571 (.A(clknet_0_net571),
    .X(clknet_1_1__leaf_net571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net575 (.A(net575),
    .X(clknet_0_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_0__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net575 (.A(clknet_0_net575),
    .X(clknet_1_1__leaf_net575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net670 (.A(net670),
    .X(clknet_0_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net670 (.A(clknet_0_net670),
    .X(clknet_1_0__leaf_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net670 (.A(clknet_0_net670),
    .X(clknet_1_1__leaf_net670));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net678 (.A(net678),
    .X(clknet_0_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_0__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_1__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net586 (.A(net586),
    .X(clknet_0_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_0__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net586 (.A(clknet_0_net586),
    .X(clknet_1_1__leaf_net586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net584 (.A(net584),
    .X(clknet_0_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net584 (.A(net757),
    .X(clknet_1_0__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net584 (.A(clknet_0_net584),
    .X(clknet_1_1__leaf_net584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net583 (.A(net583),
    .X(clknet_0_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net583 (.A(clknet_0_net583),
    .X(clknet_1_0__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net583 (.A(net759),
    .X(clknet_1_1__leaf_net583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net565 (.A(net565),
    .X(clknet_0_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_0__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_1__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net542 (.A(net542),
    .X(clknet_0_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_0__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_1__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net649 (.A(net649),
    .X(clknet_0_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_0__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net649 (.A(clknet_0_net649),
    .X(clknet_1_1__leaf_net649));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net549 (.A(net549),
    .X(clknet_0_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_0__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net549 (.A(clknet_0_net549),
    .X(clknet_1_1__leaf_net549));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net555 (.A(net555),
    .X(clknet_0_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_0__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net555 (.A(clknet_0_net555),
    .X(clknet_1_1__leaf_net555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net556 (.A(net556),
    .X(clknet_0_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_0__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net556 (.A(clknet_0_net556),
    .X(clknet_1_1__leaf_net556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net551 (.A(net551),
    .X(clknet_0_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_0__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net551 (.A(clknet_0_net551),
    .X(clknet_1_1__leaf_net551));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net548 (.A(net548),
    .X(clknet_0_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_0__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net548 (.A(clknet_0_net548),
    .X(clknet_1_1__leaf_net548));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net547 (.A(net547),
    .X(clknet_0_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_0__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net547 (.A(clknet_0_net547),
    .X(clknet_1_1__leaf_net547));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net545 (.A(net545),
    .X(clknet_0_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_0__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net545 (.A(clknet_0_net545),
    .X(clknet_1_1__leaf_net545));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net335 (.A(net335),
    .X(clknet_0_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_0__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net335 (.A(clknet_0_net335),
    .X(clknet_1_1__leaf_net335));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net336 (.A(net336),
    .X(clknet_0_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_0__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net336 (.A(clknet_0_net336),
    .X(clknet_1_1__leaf_net336));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net347 (.A(net347),
    .X(clknet_0_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_0__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net347 (.A(clknet_0_net347),
    .X(clknet_1_1__leaf_net347));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net338 (.A(net338),
    .X(clknet_0_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_0__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net338 (.A(clknet_0_net338),
    .X(clknet_1_1__leaf_net338));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net337 (.A(net337),
    .X(clknet_0_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_0__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_1__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net334 (.A(net334),
    .X(clknet_0_net334));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net334 (.A(clknet_0_net334),
    .X(clknet_1_0__leaf_net334));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net334 (.A(clknet_0_net334),
    .X(clknet_1_1__leaf_net334));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(clknet_0_net594),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(clknet_0_net584),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(clknet_0_net589),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(clknet_0_net583),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net468),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net476),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net715),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net688),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net357),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net391),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net302),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net507),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net642),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net432),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net506),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net504),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net308),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net319),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net514),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net516),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net473),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net482),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net298),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net313),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net316),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net466),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net710),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net419),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net400),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net393),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net501),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net222),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net716),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net693),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net315),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net692),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net314),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net709),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net424),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net153),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net362),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net317),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net475),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net394),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net284),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net410),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net714),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net292),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net415),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net520),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net433),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net641),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net309),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net483),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net432),
    .X(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_Q (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_SCE (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_D (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_SCD (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_X (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_DE (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_C (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_X (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_C1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_B (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A0 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_C (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_C (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_SCD (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_X (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_D_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_C1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_C_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_X (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_SCE (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_X (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_X (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_D1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_C (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_SET_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
