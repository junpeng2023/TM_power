module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire clknet_0_clk;
 wire clknet_0_net506;
 wire clknet_0_net561;
 wire clknet_0_net562;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net506;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net506;
 wire clknet_1_1__leaf_net561;
 wire clknet_1_1__leaf_net562;
 wire clknet_1_1__leaf_net563;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;

 sky130_fd_sc_hd__diode_2 ANTENNA_c100_C_N (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_D_N (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_B (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_C (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_X (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_S1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_C (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_X (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_B (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_D_N (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_C (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_C (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C_N (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_D_N (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_C (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_C (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_C_N (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_D_N (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_C (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_C (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_C_N (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_D_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_C (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_C (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_C_N (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_D_N (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_D_N (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_C_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_C (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A0 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_C_N (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_C_N (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_X (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_C (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_C (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_X (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_D_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_B1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_X (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_C (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_C (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_C (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_C (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_C (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_C (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_C (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_B (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_D1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_C1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_D1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_X (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_C1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_D1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_C (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_C (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_C1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_D1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_C (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A3 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_C1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_D1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_C (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_C (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_C (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_C (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A2 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_X (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_C (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_C (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_D1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_C1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_C_N (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_D1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_C_N (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_C (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_C (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_C (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_B (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_C (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_C_N (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D_N (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_X (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_C (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_C (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_B (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_C (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_C1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_C (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_C1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_D1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_C (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_C (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_C (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_X (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_C (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_C (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_C (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_C (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_X (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_C1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_D1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_C (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_C (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_C (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_X (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_X (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_D1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_C (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_X (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_B (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_B (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_C (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_C (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_C (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_C (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_D_N (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_C (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_C (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_C (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_C_N (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_D_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_C (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_C (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_C_N (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_D_N (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_C (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_C (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_D_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_X (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_C1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_B1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_C1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_C1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_D1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_C1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_D1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_D1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_C_N (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_D_N (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_RESET_B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_SCD (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_B (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_C_N (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_X (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_C (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_C1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_D1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_C1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_D1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_C1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_CLK_N (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_D (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_RESET_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SCD (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SCE (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SET_B (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_RESET_B (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_SCD (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_C_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_D_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_C_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_C (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_B (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_X (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_B (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_D_N (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_C (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_B (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_C (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_C (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_C_N (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_D_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_C (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_C (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_C (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_C (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_C_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_D_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_C (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_B (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_C_N (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_D_N (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_C1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_SCD (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_D_N (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D_N (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_C_N (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_D_N (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_B (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_D_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_C_N (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_B (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_C_N (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_D_N (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_C1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_C1 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_B (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_D_N (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCD (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCE (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A3 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A3 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone10_X (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold25_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold27_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_X (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_X (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_X (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_X (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_X (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_X (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_X (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_X (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_X (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_X (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_X (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_C1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A3 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_X (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_D_N (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_S1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_SCD (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A3 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_Q_N (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_D (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_Q (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_GATE_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_GATE_N (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_GATE (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_s818_CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s819_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_Q (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_s821_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s821_Q (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_s822_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s823_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s824_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s825_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s826_GATE_N (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s827_GATE_N (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__or4bb_2 c100 (.A(net662),
    .B(net608),
    .C_N(net1034),
    .D_N(net660),
    .X(net688));
 sky130_fd_sc_hd__and2_1 c101 (.A(net629),
    .B(net648),
    .X(net699));
 sky130_fd_sc_hd__and3_4 c102 (.A(net604),
    .B(net659),
    .C(net1061),
    .X(net735));
 sky130_fd_sc_hd__and2_0 c103 (.A(net615),
    .B(net658),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c104 (.A0(net657),
    .A1(net1040),
    .A2(net605),
    .A3(net615),
    .S0(net659),
    .S1(net1033),
    .X(net1));
 sky130_fd_sc_hd__and3_1 c105 (.A(net1041),
    .B(net1050),
    .C(net1047),
    .X(net2));
 sky130_fd_sc_hd__and2_1 c106 (.A(net735),
    .B(net601),
    .X(net3));
 sky130_fd_sc_hd__and2_0 c107 (.A(net664),
    .B(net735),
    .X(net703));
 sky130_fd_sc_hd__and2_1 c108 (.A(net1),
    .B(net607),
    .X(net728));
 sky130_fd_sc_hd__mux4_2 c109 (.A0(net631),
    .A1(net653),
    .A2(net2),
    .A3(net728),
    .S0(net663),
    .S1(net1041),
    .X(net722));
 sky130_fd_sc_hd__and2_0 c110 (.A(net1055),
    .B(net603),
    .X(net704));
 sky130_fd_sc_hd__and2_0 c111 (.A(net657),
    .B(net623),
    .X(net4));
 sky130_fd_sc_hd__and2_0 c112 (.A(net1062),
    .B(net1039),
    .X(net721));
 sky130_fd_sc_hd__and2_0 c113 (.A(net595),
    .B(net623),
    .X(net5));
 sky130_fd_sc_hd__and2_0 c114 (.A(net587),
    .B(net722),
    .X(net701));
 sky130_fd_sc_hd__and2_0 c115 (.A(net4),
    .B(net620),
    .X(net6));
 sky130_fd_sc_hd__and2_0 c116 (.A(net571),
    .B(net703),
    .X(net7));
 sky130_fd_sc_hd__and2_0 c117 (.A(net648),
    .B(net605),
    .X(net736));
 sky130_fd_sc_hd__and2_1 c118 (.A(net662),
    .B(net5),
    .X(net731));
 sky130_fd_sc_hd__and2_1 c119 (.A(net731),
    .B(net645),
    .X(net8));
 sky130_fd_sc_hd__and2_1 c120 (.A(net8),
    .B(net648),
    .X(net695));
 sky130_fd_sc_hd__and2_0 c121 (.A(net1),
    .B(net8),
    .X(net9));
 sky130_fd_sc_hd__and2_0 c122 (.A(net620),
    .B(net8),
    .X(net10));
 sky130_fd_sc_hd__and2_0 c123 (.A(net9),
    .B(net605),
    .X(net710));
 sky130_fd_sc_hd__and2_0 c124 (.A(net9),
    .B(net10),
    .X(net717));
 sky130_fd_sc_hd__and2_0 c125 (.A(net10),
    .B(net595),
    .X(net11));
 sky130_fd_sc_hd__and2_0 c126 (.A(net6),
    .B(net8),
    .X(net715));
 sky130_fd_sc_hd__and2_1 c127 (.A(net5),
    .B(net1041),
    .X(net693));
 sky130_fd_sc_hd__and3_1 c128 (.A(net2),
    .B(net693),
    .C(net717),
    .X(net737));
 sky130_fd_sc_hd__and2_1 c129 (.A(net7),
    .B(net737),
    .X(net730));
 sky130_fd_sc_hd__and2_0 c130 (.A(net11),
    .B(net10),
    .X(net12));
 sky130_fd_sc_hd__and3_1 c131 (.A(net12),
    .B(net603),
    .C(net737),
    .X(net712));
 sky130_fd_sc_hd__and2_1 c132 (.A(net633),
    .B(net1043),
    .X(net13));
 sky130_fd_sc_hd__and2_4 c133 (.A(net1057),
    .B(net1060),
    .X(net738));
 sky130_fd_sc_hd__and2_4 c134 (.A(net738),
    .B(net1047),
    .X(net14));
 sky130_fd_sc_hd__and2_1 c135 (.A(net600),
    .B(net1056),
    .X(net15));
 sky130_fd_sc_hd__and2_4 c136 (.A(net14),
    .B(net738),
    .X(net16));
 sky130_fd_sc_hd__and2_1 c137 (.A(net1038),
    .B(net1044),
    .X(net17));
 sky130_fd_sc_hd__and3_1 c138 (.A(net16),
    .B(net1031),
    .C(net1049),
    .X(net18));
 sky130_fd_sc_hd__and2_1 c139 (.A(net13),
    .B(net570),
    .X(net19));
 sky130_fd_sc_hd__and2_1 c140 (.A(net1066),
    .B(net14),
    .X(net729));
 sky130_fd_sc_hd__and2_1 c141 (.A(net570),
    .B(net14),
    .X(net732));
 sky130_fd_sc_hd__or4bb_1 c142 (.A(net1037),
    .B(net1047),
    .C_N(net13),
    .D_N(net729),
    .X(net20));
 sky130_fd_sc_hd__and2_1 c143 (.A(net1043),
    .B(net1020),
    .X(net21));
 sky130_fd_sc_hd__and3_1 c144 (.A(net577),
    .B(net573),
    .C(net1011),
    .X(net22));
 sky130_fd_sc_hd__and2_1 c145 (.A(net577),
    .B(net16),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net1030),
    .A1(net1067),
    .A2(net1021),
    .A3(net1046),
    .S0(net1037),
    .S1(net14),
    .X(net24));
 sky130_fd_sc_hd__and2_1 c147 (.A(net1014),
    .B(net729),
    .X(net25));
 sky130_fd_sc_hd__and2_4 c148 (.A(net729),
    .B(net1010),
    .X(net26));
 sky130_fd_sc_hd__and3_2 c149 (.A(net25),
    .B(net24),
    .C(net1010),
    .X(net27));
 sky130_fd_sc_hd__or4bb_4 c150 (.A(net22),
    .B(net25),
    .C_N(net1020),
    .D_N(net1010),
    .X(net685));
 sky130_fd_sc_hd__and3_1 c151 (.A(net24),
    .B(net1000),
    .C(net1010),
    .X(net28));
 sky130_fd_sc_hd__and3_1 c152 (.A(net25),
    .B(net1046),
    .C(net1021),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net994),
    .A1(net24),
    .A2(net22),
    .A3(net27),
    .S0(net999),
    .S1(net26),
    .X(net682));
 sky130_fd_sc_hd__and2_1 c154 (.A(net603),
    .B(net1061),
    .X(net30));
 sky130_fd_sc_hd__and2_1 c155 (.A(net593),
    .B(net577),
    .X(net733));
 sky130_fd_sc_hd__and2_1 c156 (.A(net577),
    .B(net1065),
    .X(net31));
 sky130_fd_sc_hd__or4bb_4 c157 (.A(net582),
    .B(net1047),
    .C_N(net597),
    .D_N(net1025),
    .X(net32));
 sky130_fd_sc_hd__and2_4 c158 (.A(net32),
    .B(net594),
    .X(net724));
 sky130_fd_sc_hd__and2_1 c159 (.A(net13),
    .B(net1025),
    .X(net33));
 sky130_fd_sc_hd__and2_1 c160 (.A(net1044),
    .B(net767),
    .X(net34));
 sky130_fd_sc_hd__and2_0 c161 (.A(net1054),
    .B(net1061),
    .X(net35));
 sky130_fd_sc_hd__and2_2 c162 (.A(net35),
    .B(net33),
    .X(net36));
 sky130_fd_sc_hd__and2_1 c163 (.A(net733),
    .B(net519),
    .X(net37));
 sky130_fd_sc_hd__and2_1 c164 (.A(net584),
    .B(net583),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net724),
    .A1(net37),
    .A2(net31),
    .A3(net26),
    .S0(net1025),
    .S1(net1055),
    .X(net39));
 sky130_fd_sc_hd__and3_1 c166 (.A(net32),
    .B(net604),
    .C(net1025),
    .X(net40));
 sky130_fd_sc_hd__or4bb_1 c167 (.A(net38),
    .B(net33),
    .C_N(net767),
    .D_N(net30),
    .X(net41));
 sky130_fd_sc_hd__and2_1 c168 (.A(net579),
    .B(net733),
    .X(net713));
 sky130_fd_sc_hd__and3_1 c169 (.A(net30),
    .B(net604),
    .C(net41),
    .X(net42));
 sky130_fd_sc_hd__and3_4 c170 (.A(net39),
    .B(net37),
    .C(net1006),
    .X(net43));
 sky130_fd_sc_hd__and3_1 c171 (.A(net30),
    .B(net41),
    .C(net1005),
    .X(net44));
 sky130_fd_sc_hd__and3_4 c172 (.A(net993),
    .B(net594),
    .C(net31),
    .X(net45));
 sky130_fd_sc_hd__or4bb_2 c173 (.A(net45),
    .B(net1063),
    .C_N(net593),
    .D_N(net998),
    .X(net46));
 sky130_fd_sc_hd__and3_1 c174 (.A(net45),
    .B(net1008),
    .C(net39),
    .X(net734));
 sky130_fd_sc_hd__and3_1 c175 (.A(net734),
    .B(net45),
    .C(net46),
    .X(net47));
 sky130_fd_sc_hd__and2_1 c176 (.A(net24),
    .B(net620),
    .X(net48));
 sky130_fd_sc_hd__and2_4 c177 (.A(net734),
    .B(net633),
    .X(net49));
 sky130_fd_sc_hd__and3_2 c178 (.A(net620),
    .B(net627),
    .C(net998),
    .X(net50));
 sky130_fd_sc_hd__and2_0 c179 (.A(net600),
    .B(net628),
    .X(net51));
 sky130_fd_sc_hd__and3_1 c180 (.A(net625),
    .B(net18),
    .C(net39),
    .X(net52));
 sky130_fd_sc_hd__and2_2 c181 (.A(net51),
    .B(net624),
    .X(net673));
 sky130_fd_sc_hd__and2_1 c182 (.A(net614),
    .B(net673),
    .X(net53));
 sky130_fd_sc_hd__and2_1 c183 (.A(net52),
    .B(net614),
    .X(net54));
 sky130_fd_sc_hd__and2_4 c184 (.A(net49),
    .B(net22),
    .X(net55));
 sky130_fd_sc_hd__and3_2 c185 (.A(net1037),
    .B(net625),
    .C(net583),
    .X(net726));
 sky130_fd_sc_hd__and3_1 c186 (.A(net54),
    .B(net49),
    .C(net53),
    .X(net56));
 sky130_fd_sc_hd__and3_1 c187 (.A(net26),
    .B(net53),
    .C(net726),
    .X(net57));
 sky130_fd_sc_hd__and2_2 c188 (.A(net53),
    .B(net1065),
    .X(net58));
 sky130_fd_sc_hd__or4bb_4 c189 (.A(net22),
    .B(net55),
    .C_N(net996),
    .D_N(net1054),
    .X(net59));
 sky130_fd_sc_hd__and3_1 c190 (.A(net619),
    .B(net615),
    .C(net1027),
    .X(net60));
 sky130_fd_sc_hd__and2_1 c191 (.A(net56),
    .B(net993),
    .X(net61));
 sky130_fd_sc_hd__and3_1 c192 (.A(net726),
    .B(net50),
    .C(net767),
    .X(net62));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net38),
    .A1(net61),
    .A2(net606),
    .A3(net1065),
    .S0(net59),
    .S1(net767),
    .X(net63));
 sky130_fd_sc_hd__and3_1 c194 (.A(net624),
    .B(net53),
    .C(net996),
    .X(net64));
 sky130_fd_sc_hd__and3_1 c195 (.A(net60),
    .B(net754),
    .C(net38),
    .X(net65));
 sky130_fd_sc_hd__or4bb_4 c196 (.A(net996),
    .B(net63),
    .C_N(net65),
    .D_N(net1052),
    .X(net66));
 sky130_fd_sc_hd__or4bb_4 c197 (.A(net1028),
    .B(net66),
    .C_N(net64),
    .D_N(net59),
    .X(net67));
 sky130_fd_sc_hd__and2_2 c198 (.A(net639),
    .B(net1068),
    .X(net709));
 sky130_fd_sc_hd__and2_1 c199 (.A(net630),
    .B(net50),
    .X(net708));
 sky130_fd_sc_hd__and2_0 c200 (.A(net635),
    .B(net709),
    .X(net68));
 sky130_fd_sc_hd__and3_1 c201 (.A(net993),
    .B(net611),
    .C(net709),
    .X(net711));
 sky130_fd_sc_hd__and2_0 c202 (.A(net65),
    .B(net711),
    .X(net69));
 sky130_fd_sc_hd__and2_0 c203 (.A(net61),
    .B(net58),
    .X(net70));
 sky130_fd_sc_hd__and2_1 c204 (.A(net638),
    .B(net637),
    .X(net71));
 sky130_fd_sc_hd__and2_0 c205 (.A(net35),
    .B(net724),
    .X(net72));
 sky130_fd_sc_hd__and2_1 c206 (.A(net69),
    .B(net709),
    .X(net73));
 sky130_fd_sc_hd__and2_1 c207 (.A(net47),
    .B(net53),
    .X(net74));
 sky130_fd_sc_hd__and3_1 c208 (.A(net70),
    .B(net636),
    .C(net1065),
    .X(net75));
 sky130_fd_sc_hd__and2_1 c209 (.A(net581),
    .B(net69),
    .X(net76));
 sky130_fd_sc_hd__and2_0 c210 (.A(net73),
    .B(net75),
    .X(net77));
 sky130_fd_sc_hd__and2_1 c211 (.A(net958),
    .B(net635),
    .X(net706));
 sky130_fd_sc_hd__and2_0 c212 (.A(net77),
    .B(net649),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net74),
    .A1(net78),
    .A2(net70),
    .A3(net1027),
    .S0(net958),
    .S1(net73),
    .X(net79));
 sky130_fd_sc_hd__mux4_2 c214 (.A0(net628),
    .A1(net708),
    .A2(net991),
    .A3(net71),
    .S0(net650),
    .S1(net76),
    .X(net698));
 sky130_fd_sc_hd__and2_1 c215 (.A(net71),
    .B(net955),
    .X(net80));
 sky130_fd_sc_hd__and2_1 c216 (.A(net72),
    .B(net651),
    .X(net81));
 sky130_fd_sc_hd__and2_1 c217 (.A(net81),
    .B(net711),
    .X(net82));
 sky130_fd_sc_hd__and3_1 c218 (.A(net79),
    .B(net82),
    .C(net81),
    .X(net83));
 sky130_fd_sc_hd__and3_2 c219 (.A(net82),
    .B(net83),
    .C(net81),
    .X(net84));
 sky130_fd_sc_hd__or4bb_1 c220 (.A(net39),
    .B(net74),
    .C_N(net659),
    .D_N(net656),
    .X(net725));
 sky130_fd_sc_hd__or4bb_1 c221 (.A(net653),
    .B(net68),
    .C_N(net735),
    .D_N(net1071),
    .X(net85));
 sky130_fd_sc_hd__and2_1 c222 (.A(net68),
    .B(net595),
    .X(net86));
 sky130_fd_sc_hd__and3_1 c223 (.A(net634),
    .B(net1040),
    .C(net1065),
    .X(net87));
 sky130_fd_sc_hd__and2_0 c224 (.A(net86),
    .B(net1040),
    .X(net88));
 sky130_fd_sc_hd__and2_0 c225 (.A(net1012),
    .B(net660),
    .X(net89));
 sky130_fd_sc_hd__and2_2 c226 (.A(net82),
    .B(net86),
    .X(net669));
 sky130_fd_sc_hd__and2_0 c227 (.A(net87),
    .B(net1029),
    .X(net90));
 sky130_fd_sc_hd__and2_1 c228 (.A(net608),
    .B(net86),
    .X(net91));
 sky130_fd_sc_hd__and3_2 c229 (.A(net90),
    .B(net85),
    .C(net991),
    .X(net702));
 sky130_fd_sc_hd__and2_1 c230 (.A(net86),
    .B(net88),
    .X(net700));
 sky130_fd_sc_hd__and2_1 c231 (.A(net85),
    .B(net700),
    .X(net92));
 sky130_fd_sc_hd__and3_2 c232 (.A(net606),
    .B(net47),
    .C(net1000),
    .X(net696));
 sky130_fd_sc_hd__and2_0 c233 (.A(net1068),
    .B(net669),
    .X(net93));
 sky130_fd_sc_hd__and2_1 c234 (.A(net51),
    .B(net606),
    .X(net94));
 sky130_fd_sc_hd__and2_1 c235 (.A(net659),
    .B(net576),
    .X(net95));
 sky130_fd_sc_hd__and3_1 c236 (.A(net748),
    .B(net95),
    .C(net608),
    .X(net723));
 sky130_fd_sc_hd__and2_1 c237 (.A(net91),
    .B(net88),
    .X(net96));
 sky130_fd_sc_hd__and2_1 c238 (.A(net91),
    .B(net92),
    .X(net727));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net999),
    .A1(net92),
    .A2(net727),
    .A3(net80),
    .S0(net964),
    .S1(net89),
    .X(net97));
 sky130_fd_sc_hd__and3_1 c240 (.A(net97),
    .B(net80),
    .C(net726),
    .X(net718));
 sky130_fd_sc_hd__or4bb_1 c241 (.A(net92),
    .B(net86),
    .C_N(net718),
    .D_N(net94),
    .X(net739));
 sky130_fd_sc_hd__and2_1 c264 (.A(net573),
    .B(net570),
    .X(net98));
 sky130_fd_sc_hd__and2_1 c265 (.A(net579),
    .B(net98),
    .X(net99));
 sky130_fd_sc_hd__and2_1 c266 (.A(net572),
    .B(net1063),
    .X(net719));
 sky130_fd_sc_hd__and3_1 c267 (.A(net1043),
    .B(net1049),
    .C(net98),
    .X(net697));
 sky130_fd_sc_hd__and2_2 c268 (.A(net572),
    .B(net18),
    .X(net100));
 sky130_fd_sc_hd__and2_1 c269 (.A(net98),
    .B(net1010),
    .X(net101));
 sky130_fd_sc_hd__and2_1 c270 (.A(net26),
    .B(net13),
    .X(net102));
 sky130_fd_sc_hd__and2_1 c271 (.A(net719),
    .B(net98),
    .X(net103));
 sky130_fd_sc_hd__and2_1 c272 (.A(net1042),
    .B(net1044),
    .X(net104));
 sky130_fd_sc_hd__and2_2 c273 (.A(net102),
    .B(net98),
    .X(net105));
 sky130_fd_sc_hd__and2_2 c274 (.A(net719),
    .B(net103),
    .X(net106));
 sky130_fd_sc_hd__and2_1 c275 (.A(net1036),
    .B(net102),
    .X(net107));
 sky130_fd_sc_hd__and2_1 c276 (.A(net1026),
    .B(net1038),
    .X(net108));
 sky130_fd_sc_hd__and2_1 c277 (.A(net100),
    .B(net107),
    .X(net109));
 sky130_fd_sc_hd__and2_1 c278 (.A(net105),
    .B(net1035),
    .X(net110));
 sky130_fd_sc_hd__and2_1 c279 (.A(net107),
    .B(net1036),
    .X(net111));
 sky130_fd_sc_hd__and3_1 c280 (.A(net101),
    .B(net105),
    .C(net111),
    .X(net112));
 sky130_fd_sc_hd__and2_2 c281 (.A(net1045),
    .B(net111),
    .X(net113));
 sky130_fd_sc_hd__and2_1 c282 (.A(net103),
    .B(net99),
    .X(net114));
 sky130_fd_sc_hd__and2_2 c283 (.A(net103),
    .B(net109),
    .X(net115));
 sky130_fd_sc_hd__and3_1 c284 (.A(net109),
    .B(net1036),
    .C(net990),
    .X(net116));
 sky130_fd_sc_hd__a2111o_4 c285 (.A1(net985),
    .A2(net990),
    .B1(net987),
    .C1(net1030),
    .D1(net107),
    .X(net117));
 sky130_fd_sc_hd__and2_0 c286 (.A(net519),
    .B(net45),
    .X(net118));
 sky130_fd_sc_hd__and2_2 c287 (.A(net1025),
    .B(net31),
    .X(net689));
 sky130_fd_sc_hd__and2_2 c288 (.A(net118),
    .B(net689),
    .X(net119));
 sky130_fd_sc_hd__and2_2 c289 (.A(net33),
    .B(net41),
    .X(net120));
 sky130_fd_sc_hd__and2_1 c290 (.A(net601),
    .B(net102),
    .X(net121));
 sky130_fd_sc_hd__and2_2 c291 (.A(net31),
    .B(net26),
    .X(net122));
 sky130_fd_sc_hd__and2_1 c292 (.A(net980),
    .B(net599),
    .X(net123));
 sky130_fd_sc_hd__and3_1 c293 (.A(net118),
    .B(net579),
    .C(net1061),
    .X(net124));
 sky130_fd_sc_hd__and2_1 c294 (.A(net599),
    .B(net105),
    .X(net125));
 sky130_fd_sc_hd__and2_1 c295 (.A(net121),
    .B(net33),
    .X(net126));
 sky130_fd_sc_hd__and3_1 c296 (.A(net122),
    .B(net988),
    .C(net981),
    .X(net127));
 sky130_fd_sc_hd__and3_1 c297 (.A(net37),
    .B(net33),
    .C(net738),
    .X(net128));
 sky130_fd_sc_hd__and2_1 c298 (.A(net102),
    .B(net46),
    .X(net129));
 sky130_fd_sc_hd__and3_1 c299 (.A(net41),
    .B(net586),
    .C(net1004),
    .X(net130));
 sky130_fd_sc_hd__or4bb_1 c300 (.A(net128),
    .B(net584),
    .C_N(net1036),
    .D_N(net981),
    .X(net131));
 sky130_fd_sc_hd__and2_1 c301 (.A(net1004),
    .B(net18),
    .X(net132));
 sky130_fd_sc_hd__and3_1 c302 (.A(net995),
    .B(net593),
    .C(net582),
    .X(net133));
 sky130_fd_sc_hd__and2_1 c303 (.A(net127),
    .B(net120),
    .X(net134));
 sky130_fd_sc_hd__and3_1 c304 (.A(net124),
    .B(net988),
    .C(net984),
    .X(net135));
 sky130_fd_sc_hd__and2_1 c305 (.A(net135),
    .B(net133),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net130),
    .A1(net136),
    .A2(net134),
    .A3(net995),
    .S0(net984),
    .S1(net981),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net27),
    .A1(net125),
    .A2(net995),
    .A3(net981),
    .S0(net1004),
    .S1(net767),
    .X(net138));
 sky130_fd_sc_hd__and2_2 c308 (.A(net768),
    .B(net613),
    .X(net139));
 sky130_fd_sc_hd__and3_1 c309 (.A(net52),
    .B(net578),
    .C(net1032),
    .X(net140));
 sky130_fd_sc_hd__and2_0 c310 (.A(net120),
    .B(net1050),
    .X(net141));
 sky130_fd_sc_hd__and2_4 c311 (.A(net67),
    .B(net140),
    .X(net142));
 sky130_fd_sc_hd__and2_0 c312 (.A(net627),
    .B(net623),
    .X(net143));
 sky130_fd_sc_hd__and2_1 c313 (.A(net143),
    .B(net113),
    .X(net144));
 sky130_fd_sc_hd__and2_0 c314 (.A(net609),
    .B(net142),
    .X(net145));
 sky130_fd_sc_hd__and3_1 c315 (.A(net138),
    .B(net609),
    .C(net139),
    .X(net146));
 sky130_fd_sc_hd__and2_1 c316 (.A(net49),
    .B(net143),
    .X(net147));
 sky130_fd_sc_hd__and2_0 c317 (.A(net67),
    .B(net56),
    .X(net148));
 sky130_fd_sc_hd__and2_1 c318 (.A(net55),
    .B(net1058),
    .X(net149));
 sky130_fd_sc_hd__and3_1 c319 (.A(net599),
    .B(net148),
    .C(net988),
    .X(net150));
 sky130_fd_sc_hd__and3_2 c320 (.A(net139),
    .B(net623),
    .C(net1028),
    .X(net151));
 sky130_fd_sc_hd__and3_1 c321 (.A(net142),
    .B(net607),
    .C(net673),
    .X(net152));
 sky130_fd_sc_hd__and2_0 c322 (.A(net1063),
    .B(net151),
    .X(net153));
 sky130_fd_sc_hd__and2_0 c323 (.A(net109),
    .B(net16),
    .X(net154));
 sky130_fd_sc_hd__and3_1 c324 (.A(net18),
    .B(net1005),
    .C(net982),
    .X(net155));
 sky130_fd_sc_hd__and2_1 c325 (.A(net602),
    .B(net984),
    .X(net156));
 sky130_fd_sc_hd__and2_0 c326 (.A(net975),
    .B(net140),
    .X(net707));
 sky130_fd_sc_hd__and3_1 c327 (.A(net151),
    .B(net961),
    .C(net152),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net156),
    .A1(net149),
    .A2(net1062),
    .A3(net599),
    .S0(net139),
    .S1(net621),
    .X(net158));
 sky130_fd_sc_hd__and3_1 c329 (.A(net141),
    .B(net158),
    .C(net151),
    .X(net159));
 sky130_fd_sc_hd__and2_1 c330 (.A(net54),
    .B(net955),
    .X(net160));
 sky130_fd_sc_hd__and2_0 c331 (.A(net79),
    .B(net156),
    .X(net161));
 sky130_fd_sc_hd__a2111o_2 c332 (.A1(net83),
    .A2(net1074),
    .B1(net1028),
    .C1(net56),
    .D1(net1079),
    .X(net162));
 sky130_fd_sc_hd__and3_1 c333 (.A(net53),
    .B(net61),
    .C(net982),
    .X(net163));
 sky130_fd_sc_hd__a2111o_2 c334 (.A1(net583),
    .A2(net83),
    .B1(net980),
    .C1(net1080),
    .D1(net960),
    .X(net687));
 sky130_fd_sc_hd__a2111o_1 c335 (.A1(net48),
    .A2(net139),
    .B1(net123),
    .C1(net144),
    .D1(net119),
    .X(net164));
 sky130_fd_sc_hd__and2_1 c336 (.A(net610),
    .B(net73),
    .X(net165));
 sky130_fd_sc_hd__and3_1 c337 (.A(net156),
    .B(net993),
    .C(net161),
    .X(net166));
 sky130_fd_sc_hd__a2111o_1 c338 (.A1(net107),
    .A2(net982),
    .B1(net992),
    .C1(net58),
    .D1(net981),
    .X(net667));
 sky130_fd_sc_hd__and3_1 c339 (.A(net149),
    .B(net27),
    .C(net687),
    .X(net167));
 sky130_fd_sc_hd__and3_1 c340 (.A(net157),
    .B(net151),
    .C(net961),
    .X(net168));
 sky130_fd_sc_hd__and2_1 c341 (.A(net27),
    .B(net966),
    .X(net169));
 sky130_fd_sc_hd__and3_1 c342 (.A(net637),
    .B(net749),
    .C(net966),
    .X(net170));
 sky130_fd_sc_hd__and3_1 c343 (.A(net113),
    .B(net165),
    .C(net966),
    .X(net171));
 sky130_fd_sc_hd__and3_2 c344 (.A(net160),
    .B(net169),
    .C(net641),
    .X(net172));
 sky130_fd_sc_hd__a2111o_2 c345 (.A1(net144),
    .A2(net146),
    .B1(net626),
    .C1(net966),
    .D1(net960),
    .X(net173));
 sky130_fd_sc_hd__and3_1 c346 (.A(net75),
    .B(net165),
    .C(net171),
    .X(net174));
 sky130_fd_sc_hd__and3_1 c347 (.A(net174),
    .B(net160),
    .C(net687),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c348 (.A(net161),
    .B(net48),
    .C(net966),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_1 c349 (.A(net1024),
    .X(net176));
 sky130_fd_sc_hd__buf_1 c350 (.A(net1024),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net171),
    .A1(net713),
    .A2(net177),
    .A3(net966),
    .S0(net172),
    .S1(net119),
    .X(net178));
 sky130_fd_sc_hd__a2111o_1 c352 (.A1(net93),
    .A2(net640),
    .B1(net722),
    .C1(net642),
    .D1(net696),
    .X(net179));
 sky130_fd_sc_hd__and3_1 c353 (.A(net134),
    .B(net720),
    .C(net966),
    .X(net180));
 sky130_fd_sc_hd__and3_1 c354 (.A(net168),
    .B(net632),
    .C(net955),
    .X(net181));
 sky130_fd_sc_hd__and3_1 c355 (.A(net179),
    .B(net151),
    .C(net956),
    .X(net182));
 sky130_fd_sc_hd__and2_0 c356 (.A(net621),
    .B(net626),
    .X(net183));
 sky130_fd_sc_hd__and3_1 c357 (.A(net56),
    .B(net43),
    .C(net173),
    .X(net684));
 sky130_fd_sc_hd__mux4_2 c358 (.A0(net0),
    .A1(net999),
    .A2(net650),
    .A3(net1067),
    .S0(net574),
    .S1(net1040),
    .X(net184));
 sky130_fd_sc_hd__and3_1 c359 (.A(net654),
    .B(net127),
    .C(net184),
    .X(net185));
 sky130_fd_sc_hd__and3_1 c360 (.A(net756),
    .B(net621),
    .C(net642),
    .X(net186));
 sky130_fd_sc_hd__and3_1 c361 (.A(net117),
    .B(net654),
    .C(net183),
    .X(net187));
 sky130_fd_sc_hd__mux4_2 c362 (.A0(net88),
    .A1(net575),
    .A2(net85),
    .A3(net980),
    .S0(net702),
    .S1(net1034),
    .X(net188));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net146),
    .A1(net1072),
    .A2(net1079),
    .A3(net650),
    .S0(net991),
    .S1(net80),
    .X(net705));
 sky130_fd_sc_hd__a2111o_4 c364 (.A1(net184),
    .A2(net168),
    .B1(net966),
    .C1(net151),
    .D1(net706),
    .X(net189));
 sky130_fd_sc_hd__and3_1 c365 (.A(net89),
    .B(net183),
    .C(net94),
    .X(net691));
 sky130_fd_sc_hd__and2_0 c366 (.A(net94),
    .B(net185),
    .X(net190));
 sky130_fd_sc_hd__and3_1 c367 (.A(net166),
    .B(net1030),
    .C(net957),
    .X(net191));
 sky130_fd_sc_hd__and3_1 c368 (.A(net190),
    .B(net189),
    .C(net151),
    .X(net192));
 sky130_fd_sc_hd__and3_1 c369 (.A(net80),
    .B(net85),
    .C(net189),
    .X(net193));
 sky130_fd_sc_hd__and2_0 c370 (.A(net165),
    .B(net91),
    .X(net194));
 sky130_fd_sc_hd__buf_1 c371 (.A(net774),
    .X(net195));
 sky130_fd_sc_hd__and3_1 c372 (.A(net187),
    .B(net189),
    .C(net718),
    .X(net196));
 sky130_fd_sc_hd__a2111o_1 c373 (.A1(net1065),
    .A2(net196),
    .B1(net61),
    .C1(net195),
    .D1(net189),
    .X(net197));
 sky130_fd_sc_hd__and2_1 c396 (.A(net114),
    .B(net1068),
    .X(net198));
 sky130_fd_sc_hd__and2_1 c397 (.A(net572),
    .B(net1010),
    .X(net199));
 sky130_fd_sc_hd__and3_2 c398 (.A(net199),
    .B(net98),
    .C(net15),
    .X(net200));
 sky130_fd_sc_hd__and2_1 c399 (.A(net1045),
    .B(net985),
    .X(net201));
 sky130_fd_sc_hd__and2_2 c400 (.A(net111),
    .B(net1026),
    .X(net202));
 sky130_fd_sc_hd__and2_2 c401 (.A(net1070),
    .B(net1013),
    .X(net681));
 sky130_fd_sc_hd__and2_0 c402 (.A(net98),
    .B(net202),
    .X(net203));
 sky130_fd_sc_hd__and2_2 c403 (.A(net198),
    .B(net983),
    .X(net204));
 sky130_fd_sc_hd__and2_1 c404 (.A(net114),
    .B(net1015),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c405 (.A(net519),
    .B(net1070),
    .X(net206));
 sky130_fd_sc_hd__a2111o_2 c406 (.A1(net987),
    .A2(net114),
    .B1(net202),
    .C1(net199),
    .D1(net1003),
    .X(net207));
 sky130_fd_sc_hd__and2_2 c407 (.A(net202),
    .B(net199),
    .X(net686));
 sky130_fd_sc_hd__and2_0 c408 (.A(net200),
    .B(net202),
    .X(net208));
 sky130_fd_sc_hd__and2_1 c409 (.A(net206),
    .B(net1003),
    .X(net209));
 sky130_fd_sc_hd__and2_2 c410 (.A(net200),
    .B(net202),
    .X(net210));
 sky130_fd_sc_hd__and2_0 c411 (.A(net203),
    .B(net205),
    .X(net211));
 sky130_fd_sc_hd__and2_2 c412 (.A(net25),
    .B(net1042),
    .X(net692));
 sky130_fd_sc_hd__and2_1 c413 (.A(net209),
    .B(net1046),
    .X(net212));
 sky130_fd_sc_hd__and2_2 c414 (.A(net212),
    .B(net202),
    .X(net674));
 sky130_fd_sc_hd__and2_0 c415 (.A(net204),
    .B(net212),
    .X(net213));
 sky130_fd_sc_hd__and2_1 c416 (.A(net211),
    .B(net113),
    .X(net214));
 sky130_fd_sc_hd__a2111o_1 c417 (.A1(net983),
    .A2(net101),
    .B1(net692),
    .C1(net200),
    .D1(net202),
    .X(net215));
 sky130_fd_sc_hd__and2_2 c418 (.A(net995),
    .B(net1020),
    .X(net216));
 sky130_fd_sc_hd__and2_1 c419 (.A(net15),
    .B(net204),
    .X(net217));
 sky130_fd_sc_hd__and2_0 c420 (.A(net18),
    .B(net1036),
    .X(net218));
 sky130_fd_sc_hd__or4bb_1 c421 (.A(net1015),
    .B(net217),
    .C_N(net1026),
    .D_N(net978),
    .X(net219));
 sky130_fd_sc_hd__a2111o_1 c422 (.A1(net111),
    .A2(net210),
    .B1(net1014),
    .C1(net212),
    .D1(net1017),
    .X(net220));
 sky130_fd_sc_hd__and2_1 c423 (.A(net127),
    .B(net30),
    .X(net221));
 sky130_fd_sc_hd__and2_1 c424 (.A(net216),
    .B(net131),
    .X(net222));
 sky130_fd_sc_hd__and3_2 c425 (.A(net1054),
    .B(net207),
    .C(net221),
    .X(net679));
 sky130_fd_sc_hd__or4bb_2 c426 (.A(net99),
    .B(net46),
    .C_N(net679),
    .D_N(net978),
    .X(net223));
 sky130_fd_sc_hd__and3_2 c427 (.A(net973),
    .B(net218),
    .C(net121),
    .X(net224));
 sky130_fd_sc_hd__and2_1 c428 (.A(net46),
    .B(net220),
    .X(net225));
 sky130_fd_sc_hd__and2_4 c429 (.A(net219),
    .B(net220),
    .X(net226));
 sky130_fd_sc_hd__and3_1 c430 (.A(net124),
    .B(net222),
    .C(net1015),
    .X(net227));
 sky130_fd_sc_hd__and3_1 c431 (.A(net223),
    .B(net204),
    .C(net970),
    .X(net228));
 sky130_fd_sc_hd__and3_1 c432 (.A(net128),
    .B(net228),
    .C(net689),
    .X(net229));
 sky130_fd_sc_hd__mux4_2 c433 (.A0(net224),
    .A1(net970),
    .A2(net973),
    .A3(net1062),
    .S0(net1045),
    .S1(net206),
    .X(net230));
 sky130_fd_sc_hd__and2_1 c434 (.A(net225),
    .B(net124),
    .X(net231));
 sky130_fd_sc_hd__and2_1 c435 (.A(net973),
    .B(net231),
    .X(net232));
 sky130_fd_sc_hd__and2_1 c436 (.A(net232),
    .B(net132),
    .X(net233));
 sky130_fd_sc_hd__and2_0 c437 (.A(net230),
    .B(net227),
    .X(net234));
 sky130_fd_sc_hd__and2_0 c438 (.A(net229),
    .B(net234),
    .X(net235));
 sky130_fd_sc_hd__and2_1 c439 (.A(net226),
    .B(net679),
    .X(net236));
 sky130_fd_sc_hd__and2_0 c440 (.A(net1059),
    .B(net963),
    .X(net237));
 sky130_fd_sc_hd__and3_1 c441 (.A(net234),
    .B(net990),
    .C(net155),
    .X(net238));
 sky130_fd_sc_hd__and3_1 c442 (.A(net125),
    .B(net235),
    .C(net57),
    .X(net239));
 sky130_fd_sc_hd__and2_0 c443 (.A(net220),
    .B(net58),
    .X(net240));
 sky130_fd_sc_hd__and2_0 c444 (.A(net1032),
    .B(net975),
    .X(net241));
 sky130_fd_sc_hd__and3_1 c445 (.A(net159),
    .B(net985),
    .C(net982),
    .X(net242));
 sky130_fd_sc_hd__and3_1 c446 (.A(net133),
    .B(net100),
    .C(net16),
    .X(net243));
 sky130_fd_sc_hd__and2_1 c447 (.A(net148),
    .B(net222),
    .X(net244));
 sky130_fd_sc_hd__and2_2 c448 (.A(net616),
    .B(net106),
    .X(net666));
 sky130_fd_sc_hd__or4bb_1 c449 (.A(net238),
    .B(net666),
    .C_N(net42),
    .D_N(net961),
    .X(net245));
 sky130_fd_sc_hd__and2_2 c450 (.A(net240),
    .B(net230),
    .X(net675));
 sky130_fd_sc_hd__and2_1 c451 (.A(net218),
    .B(net113),
    .X(net246));
 sky130_fd_sc_hd__a2111o_1 c452 (.A1(net970),
    .A2(net152),
    .B1(net975),
    .C1(net139),
    .D1(net238),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c453 (.A(net245),
    .B(net673),
    .C(net769),
    .X(net248));
 sky130_fd_sc_hd__and3_1 c454 (.A(net247),
    .B(net963),
    .C(net220),
    .X(net249));
 sky130_fd_sc_hd__and3_1 c455 (.A(net247),
    .B(net153),
    .C(net126),
    .X(net250));
 sky130_fd_sc_hd__and2_0 c456 (.A(net249),
    .B(net1075),
    .X(net251));
 sky130_fd_sc_hd__and3_1 c457 (.A(net131),
    .B(net251),
    .C(net602),
    .X(net252));
 sky130_fd_sc_hd__and2_0 c458 (.A(net243),
    .B(net245),
    .X(net253));
 sky130_fd_sc_hd__and3_1 c459 (.A(net1042),
    .B(net15),
    .C(net246),
    .X(net254));
 sky130_fd_sc_hd__and3_4 c460 (.A(net250),
    .B(net249),
    .C(net254),
    .X(net255));
 sky130_fd_sc_hd__a2111o_4 c461 (.A1(net253),
    .A2(net1076),
    .B1(net30),
    .C1(net981),
    .D1(net751),
    .X(net256));
 sky130_fd_sc_hd__and3_1 c462 (.A(net78),
    .B(net610),
    .C(net636),
    .X(net257));
 sky130_fd_sc_hd__and2_0 c463 (.A(net251),
    .B(net139),
    .X(net258));
 sky130_fd_sc_hd__and3_1 c464 (.A(net586),
    .B(net30),
    .C(net1036),
    .X(net259));
 sky130_fd_sc_hd__and3_1 c465 (.A(net16),
    .B(net240),
    .C(net162),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net552),
    .X(net261));
 sky130_fd_sc_hd__a2111o_1 c467 (.A1(net176),
    .A2(net100),
    .B1(net647),
    .C1(net232),
    .D1(net961),
    .X(net262));
 sky130_fd_sc_hd__buf_1 c468 (.A(net680),
    .X(net263));
 sky130_fd_sc_hd__a2111o_1 c469 (.A1(net64),
    .A2(net984),
    .B1(net692),
    .C1(net1059),
    .D1(net697),
    .X(net264));
 sky130_fd_sc_hd__and3_1 c470 (.A(net209),
    .B(net168),
    .C(net753),
    .X(net265));
 sky130_fd_sc_hd__and3_2 c471 (.A(net265),
    .B(net636),
    .C(net974),
    .X(net266));
 sky130_fd_sc_hd__and3_1 c472 (.A(net259),
    .B(net263),
    .C(net139),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net248),
    .A1(net575),
    .A2(net139),
    .A3(net963),
    .S0(net239),
    .S1(net1052),
    .X(net268));
 sky130_fd_sc_hd__dlymetal6s2s_1 c474 (.A(net552),
    .X(net269));
 sky130_fd_sc_hd__and3_1 c475 (.A(net205),
    .B(net262),
    .C(net264),
    .X(net270));
 sky130_fd_sc_hd__and3_1 c476 (.A(net58),
    .B(net262),
    .C(net675),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 c477 (.A(net552),
    .X(net272));
 sky130_fd_sc_hd__and3_1 c478 (.A(net267),
    .B(net272),
    .C(net259),
    .X(net273));
 sky130_fd_sc_hd__and2_2 c479 (.A(net177),
    .B(net229),
    .X(net668));
 sky130_fd_sc_hd__and3_2 c480 (.A(net162),
    .B(net586),
    .C(net269),
    .X(net670));
 sky130_fd_sc_hd__and3_1 c481 (.A(net100),
    .B(net273),
    .C(net607),
    .X(net274));
 sky130_fd_sc_hd__and3_1 c482 (.A(net274),
    .B(net270),
    .C(net269),
    .X(net275));
 sky130_fd_sc_hd__and3_1 c483 (.A(net246),
    .B(net261),
    .C(net28),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net626),
    .A1(net601),
    .A2(net960),
    .A3(net178),
    .S0(net652),
    .S1(net980),
    .X(net694));
 sky130_fd_sc_hd__and3_1 c485 (.A(net583),
    .B(net61),
    .C(net968),
    .X(net277));
 sky130_fd_sc_hd__and2_0 c486 (.A(net244),
    .B(net189),
    .X(net278));
 sky130_fd_sc_hd__and3_4 c487 (.A(net663),
    .B(net200),
    .C(net1040),
    .X(net672));
 sky130_fd_sc_hd__and2_1 c488 (.A(net607),
    .B(net3),
    .X(net279));
 sky130_fd_sc_hd__a2111o_2 c489 (.A1(net181),
    .A2(net277),
    .B1(net96),
    .C1(net672),
    .D1(net1040),
    .X(net280));
 sky130_fd_sc_hd__and3_1 c490 (.A(net652),
    .B(net95),
    .C(net696),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 c491 (.A(net541),
    .X(net282));
 sky130_fd_sc_hd__mux4_2 c492 (.A0(net178),
    .A1(net722),
    .A2(net663),
    .A3(net123),
    .S0(net1012),
    .S1(net189),
    .X(net283));
 sky130_fd_sc_hd__and3_1 c493 (.A(net96),
    .B(net661),
    .C(net224),
    .X(net678));
 sky130_fd_sc_hd__and2_1 c494 (.A(net182),
    .B(net602),
    .X(net284));
 sky130_fd_sc_hd__and3_1 c495 (.A(net228),
    .B(net224),
    .C(net189),
    .X(net285));
 sky130_fd_sc_hd__and3_1 c496 (.A(net123),
    .B(net276),
    .C(net1062),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net627),
    .A1(net191),
    .A2(net955),
    .A3(net652),
    .S0(net633),
    .S1(net968),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net658),
    .A1(net286),
    .A2(net189),
    .A3(net955),
    .S0(net627),
    .S1(net694),
    .X(net288));
 sky130_fd_sc_hd__and2_1 c499 (.A(net95),
    .B(net92),
    .X(net289));
 sky130_fd_sc_hd__and3_1 c500 (.A(net186),
    .B(net194),
    .C(net1029),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 c501 (.A(net541),
    .X(net291));
 sky130_fd_sc_hd__and2_0 c502 (.A(net3),
    .B(net680),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 c503 (.A(net1024),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net292),
    .A1(net293),
    .A2(net173),
    .A3(net163),
    .S0(net972),
    .S1(net285),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net254),
    .A1(net647),
    .A2(net244),
    .A3(net283),
    .S0(net645),
    .S1(net688),
    .X(net295));
 sky130_fd_sc_hd__and2_1 c528 (.A(net213),
    .B(net987),
    .X(net296));
 sky130_fd_sc_hd__and2_1 c529 (.A(net203),
    .B(net211),
    .X(net297));
 sky130_fd_sc_hd__and2_1 c530 (.A(net999),
    .B(net297),
    .X(net298));
 sky130_fd_sc_hd__and2_0 c531 (.A(net1049),
    .B(net215),
    .X(net299));
 sky130_fd_sc_hd__and2_1 c532 (.A(net573),
    .B(net1011),
    .X(net300));
 sky130_fd_sc_hd__and2_0 c533 (.A(net296),
    .B(net300),
    .X(net301));
 sky130_fd_sc_hd__and2_1 c534 (.A(net579),
    .B(net298),
    .X(net302));
 sky130_fd_sc_hd__and2_1 c535 (.A(net298),
    .B(net1001),
    .X(net303));
 sky130_fd_sc_hd__and2_0 c536 (.A(net983),
    .B(net1057),
    .X(net304));
 sky130_fd_sc_hd__and2_1 c537 (.A(net301),
    .B(net208),
    .X(net305));
 sky130_fd_sc_hd__and2_1 c538 (.A(net199),
    .B(net1010),
    .X(net306));
 sky130_fd_sc_hd__and2_1 c539 (.A(net302),
    .B(net213),
    .X(net307));
 sky130_fd_sc_hd__and2_1 c540 (.A(net1066),
    .B(net306),
    .X(net308));
 sky130_fd_sc_hd__a2111o_1 c541 (.A1(net117),
    .A2(net298),
    .B1(net308),
    .C1(net302),
    .D1(net1048),
    .X(net309));
 sky130_fd_sc_hd__and2_2 c542 (.A(net962),
    .B(net299),
    .X(net310));
 sky130_fd_sc_hd__and2_0 c543 (.A(net308),
    .B(net674),
    .X(net311));
 sky130_fd_sc_hd__and3_1 c544 (.A(net308),
    .B(net305),
    .C(net962),
    .X(net312));
 sky130_fd_sc_hd__and2_0 c545 (.A(net297),
    .B(net305),
    .X(net313));
 sky130_fd_sc_hd__and2_0 c546 (.A(net304),
    .B(net313),
    .X(net314));
 sky130_fd_sc_hd__and2_1 c547 (.A(net299),
    .B(net296),
    .X(net315));
 sky130_fd_sc_hd__and2_2 c548 (.A(net312),
    .B(net311),
    .X(net677));
 sky130_fd_sc_hd__and2_1 c549 (.A(net314),
    .B(net315),
    .X(net316));
 sky130_fd_sc_hd__and2_1 c550 (.A(net1045),
    .B(net236),
    .X(net317));
 sky130_fd_sc_hd__and3_1 c551 (.A(net593),
    .B(net130),
    .C(net198),
    .X(net318));
 sky130_fd_sc_hd__and2_1 c552 (.A(net231),
    .B(net207),
    .X(net319));
 sky130_fd_sc_hd__and3_1 c553 (.A(net208),
    .B(net1018),
    .C(net317),
    .X(net320));
 sky130_fd_sc_hd__a2111o_1 c554 (.A1(net212),
    .A2(net122),
    .B1(net236),
    .C1(net978),
    .D1(net317),
    .X(net321));
 sky130_fd_sc_hd__and2_0 c555 (.A(net130),
    .B(net321),
    .X(net322));
 sky130_fd_sc_hd__and2_1 c556 (.A(net309),
    .B(net14),
    .X(net323));
 sky130_fd_sc_hd__and3_1 c557 (.A(net101),
    .B(net1007),
    .C(net208),
    .X(net324));
 sky130_fd_sc_hd__and3_1 c558 (.A(net317),
    .B(net633),
    .C(net202),
    .X(net325));
 sky130_fd_sc_hd__and2_0 c559 (.A(net597),
    .B(net318),
    .X(net326));
 sky130_fd_sc_hd__and3_1 c560 (.A(net326),
    .B(net987),
    .C(net983),
    .X(net327));
 sky130_fd_sc_hd__and3_1 c561 (.A(net323),
    .B(net322),
    .C(net644),
    .X(net328));
 sky130_fd_sc_hd__and2_0 c562 (.A(net236),
    .B(net1001),
    .X(net329));
 sky130_fd_sc_hd__and2_1 c563 (.A(net327),
    .B(net298),
    .X(net330));
 sky130_fd_sc_hd__and2_1 c564 (.A(net321),
    .B(net330),
    .X(net331));
 sky130_fd_sc_hd__and3_1 c565 (.A(net326),
    .B(net328),
    .C(net978),
    .X(net332));
 sky130_fd_sc_hd__and3_1 c566 (.A(net519),
    .B(net327),
    .C(net323),
    .X(net333));
 sky130_fd_sc_hd__and2_1 c567 (.A(net333),
    .B(net332),
    .X(net334));
 sky130_fd_sc_hd__and3_1 c568 (.A(net319),
    .B(net13),
    .C(net221),
    .X(net335));
 sky130_fd_sc_hd__and3_1 c569 (.A(net328),
    .B(net217),
    .C(net969),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net334),
    .A1(net332),
    .A2(net317),
    .A3(net329),
    .S0(net226),
    .S1(net335),
    .X(net337));
 sky130_fd_sc_hd__and3_2 c571 (.A(net336),
    .B(net597),
    .C(net335),
    .X(net676));
 sky130_fd_sc_hd__and3_1 c572 (.A(net150),
    .B(net336),
    .C(net600),
    .X(net338));
 sky130_fd_sc_hd__and2_0 c573 (.A(net310),
    .B(net618),
    .X(net339));
 sky130_fd_sc_hd__and3_2 c574 (.A(net215),
    .B(net335),
    .C(net682),
    .X(net340));
 sky130_fd_sc_hd__or4bb_1 c575 (.A(net298),
    .B(net135),
    .C_N(net150),
    .D_N(net675),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net759),
    .X(net342));
 sky130_fd_sc_hd__and3_1 c577 (.A(net198),
    .B(net340),
    .C(net155),
    .X(net343));
 sky130_fd_sc_hd__and3_1 c578 (.A(net953),
    .B(net674),
    .C(net323),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 c579 (.A(net543),
    .X(net345));
 sky130_fd_sc_hd__and3_1 c580 (.A(net318),
    .B(net1015),
    .C(net1051),
    .X(net346));
 sky130_fd_sc_hd__and3_1 c581 (.A(net129),
    .B(net117),
    .C(net685),
    .X(net347));
 sky130_fd_sc_hd__and3_1 c582 (.A(net346),
    .B(net154),
    .C(net1052),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 c583 (.A(net952),
    .X(net349));
 sky130_fd_sc_hd__and3_1 c584 (.A(net343),
    .B(net1052),
    .C(net1030),
    .X(net350));
 sky130_fd_sc_hd__or4bb_4 c585 (.A(net202),
    .B(net1011),
    .C_N(net1068),
    .D_N(net349),
    .X(net351));
 sky130_fd_sc_hd__and3_1 c586 (.A(net330),
    .B(net953),
    .C(net1049),
    .X(net352));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net1018),
    .A1(net219),
    .A2(net951),
    .A3(net301),
    .S0(net351),
    .S1(net320),
    .X(net353));
 sky130_fd_sc_hd__and2_0 c588 (.A(net618),
    .B(net319),
    .X(net354));
 sky130_fd_sc_hd__mux4_2 c589 (.A0(net988),
    .A1(net987),
    .A2(net346),
    .A3(net353),
    .S0(net325),
    .S1(net677),
    .X(net671));
 sky130_fd_sc_hd__and2_1 c590 (.A(net320),
    .B(net609),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net589),
    .A1(net155),
    .A2(net340),
    .A3(net121),
    .S0(net347),
    .S1(net990),
    .X(net356));
 sky130_fd_sc_hd__and3_1 c592 (.A(net348),
    .B(net62),
    .C(net951),
    .X(net357));
 sky130_fd_sc_hd__and3_1 c593 (.A(net62),
    .B(net355),
    .C(net951),
    .X(net358));
 sky130_fd_sc_hd__or4bb_1 c594 (.A(net264),
    .B(net259),
    .C_N(net1016),
    .D_N(net757),
    .X(net359));
 sky130_fd_sc_hd__and3_1 c595 (.A(net311),
    .B(net304),
    .C(net643),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 c596 (.A(net547),
    .X(net360));
 sky130_fd_sc_hd__and3_1 c597 (.A(net158),
    .B(net226),
    .C(net257),
    .X(net361));
 sky130_fd_sc_hd__and3_1 c598 (.A(net241),
    .B(net232),
    .C(net169),
    .X(net362));
 sky130_fd_sc_hd__and2_0 c599 (.A(net313),
    .B(net221),
    .X(net363));
 sky130_fd_sc_hd__and2_2 c600 (.A(net306),
    .B(net992),
    .X(net364));
 sky130_fd_sc_hd__and3_1 c601 (.A(net235),
    .B(net137),
    .C(net268),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 c602 (.A(net547),
    .X(net366));
 sky130_fd_sc_hd__and3_1 c603 (.A(net643),
    .B(net1065),
    .C(net766),
    .X(net367));
 sky130_fd_sc_hd__and3_1 c604 (.A(net242),
    .B(net364),
    .C(net137),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net365),
    .A1(net361),
    .A2(net668),
    .A3(net1068),
    .S0(net364),
    .S1(net1042),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 c606 (.A(net547),
    .X(net370));
 sky130_fd_sc_hd__and3_1 c607 (.A(net963),
    .B(net201),
    .C(net169),
    .X(net371));
 sky130_fd_sc_hd__and3_1 c608 (.A(net354),
    .B(net257),
    .C(net364),
    .X(net372));
 sky130_fd_sc_hd__or4bb_1 c609 (.A(net352),
    .B(net371),
    .C_N(net364),
    .D_N(net972),
    .X(net373));
 sky130_fd_sc_hd__and3_1 c610 (.A(net372),
    .B(net611),
    .C(net530),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net169),
    .A1(net685),
    .A2(net233),
    .A3(net365),
    .S0(net958),
    .S1(net974),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net366),
    .A1(net1005),
    .A2(net364),
    .A3(net57),
    .S0(net972),
    .S1(net556),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 c613 (.A(net547),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 c614 (.A(net567),
    .X(net378));
 sky130_fd_sc_hd__and3_1 c615 (.A(net239),
    .B(net376),
    .C(net557),
    .X(net379));
 sky130_fd_sc_hd__a2111o_1 c616 (.A1(net1052),
    .A2(net1032),
    .B1(net668),
    .C1(net999),
    .D1(net364),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net223),
    .A1(net374),
    .A2(net581),
    .A3(net1068),
    .S0(net646),
    .S1(net964),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 c618 (.A(net564),
    .X(net683));
 sky130_fd_sc_hd__a2111o_1 c619 (.A1(net285),
    .A2(net770),
    .B1(net961),
    .C1(net670),
    .D1(net117),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net163),
    .A1(net269),
    .A2(net275),
    .A3(net669),
    .S0(net266),
    .S1(net188),
    .X(net383));
 sky130_fd_sc_hd__a2111o_1 c621 (.A1(net339),
    .A2(net381),
    .B1(net256),
    .C1(net964),
    .D1(net223),
    .X(net384));
 sky130_fd_sc_hd__a2111o_1 c622 (.A1(net331),
    .A2(net368),
    .B1(net672),
    .C1(net670),
    .D1(net997),
    .X(net385));
 sky130_fd_sc_hd__a2111o_1 c623 (.A1(net137),
    .A2(net1008),
    .B1(net957),
    .C1(net269),
    .D1(net682),
    .X(net386));
 sky130_fd_sc_hd__or4bb_1 c624 (.A(net170),
    .B(net985),
    .C_N(net1051),
    .D_N(net986),
    .X(net387));
 sky130_fd_sc_hd__sdfbbn_1 c625 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net173),
    .RESET_B(net972),
    .SCD(net957),
    .SCE(net381),
    .SET_B(net557),
    .Q(net388));
 sky130_fd_sc_hd__or4bb_1 c626 (.A(net388),
    .B(net116),
    .C_N(net1012),
    .D_N(net546),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net340),
    .A1(net362),
    .A2(net646),
    .A3(net269),
    .S0(net961),
    .S1(net542),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 c628 (.A0(net356),
    .A1(net581),
    .A2(net1008),
    .A3(net1032),
    .S0(net368),
    .S1(net961),
    .X(net391));
 sky130_fd_sc_hd__and3_1 c629 (.A(net584),
    .B(net291),
    .C(net674),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net1012),
    .A1(net364),
    .A2(net289),
    .A3(net1052),
    .S0(net1058),
    .S1(net556),
    .X(net393));
 sky130_fd_sc_hd__a2111o_1 c631 (.A1(net655),
    .A2(net353),
    .B1(net1056),
    .C1(net170),
    .D1(net977),
    .X(net394));
 sky130_fd_sc_hd__a2111o_1 c632 (.A1(net393),
    .A2(net115),
    .B1(net390),
    .C1(net999),
    .D1(net1065),
    .X(net395));
 sky130_fd_sc_hd__a2111o_1 c633 (.A1(net750),
    .A2(net204),
    .B1(net389),
    .C1(net672),
    .D1(net392),
    .X(net396));
 sky130_fd_sc_hd__sdfbbn_1 c634 (.CLK_N(clknet_2_2__leaf_clk),
    .D(net575),
    .RESET_B(net57),
    .SCD(net1049),
    .SCE(net285),
    .SET_B(net391),
    .Q(net398),
    .Q_N(net397));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net1056),
    .A1(net395),
    .A2(net284),
    .A3(net115),
    .S0(net397),
    .S1(net755),
    .X(net399));
 sky130_fd_sc_hd__sdfrbp_1 c636 (.CLK(clknet_2_2__leaf_clk),
    .D(net278),
    .RESET_B(net676),
    .SCD(net987),
    .SCE(net775),
    .Q(net400));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net776),
    .A1(net283),
    .A2(net340),
    .A3(net399),
    .S0(net391),
    .S1(net1060),
    .X(net401));
 sky130_fd_sc_hd__and2_0 c660 (.A(net578),
    .B(net106),
    .X(net402));
 sky130_fd_sc_hd__and2_1 c661 (.A(net570),
    .B(net214),
    .X(net403));
 sky130_fd_sc_hd__and2_1 c662 (.A(net1057),
    .B(net310),
    .X(net404));
 sky130_fd_sc_hd__and2_0 c663 (.A(net214),
    .B(net1014),
    .X(net405));
 sky130_fd_sc_hd__and2_0 c664 (.A(net1010),
    .B(net214),
    .X(net406));
 sky130_fd_sc_hd__and2_1 c665 (.A(net316),
    .B(net309),
    .X(net407));
 sky130_fd_sc_hd__and2_0 c666 (.A(net303),
    .B(net1003),
    .X(net408));
 sky130_fd_sc_hd__and2_1 c667 (.A(net1020),
    .B(net1003),
    .X(net409));
 sky130_fd_sc_hd__and3_1 c668 (.A(net211),
    .B(net682),
    .C(net409),
    .X(net410));
 sky130_fd_sc_hd__and3_2 c669 (.A(net408),
    .B(net1067),
    .C(net409),
    .X(net411));
 sky130_fd_sc_hd__and2_0 c670 (.A(net402),
    .B(net316),
    .X(net412));
 sky130_fd_sc_hd__and2_1 c671 (.A(net407),
    .B(net115),
    .X(net413));
 sky130_fd_sc_hd__and3_1 c672 (.A(net409),
    .B(net309),
    .C(net407),
    .X(net414));
 sky130_fd_sc_hd__and3_1 c673 (.A(net414),
    .B(net413),
    .C(net408),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(net302),
    .A1(net303),
    .A2(net312),
    .A3(net994),
    .S0(net410),
    .S1(net316),
    .X(net416));
 sky130_fd_sc_hd__and2_0 c675 (.A(net410),
    .B(net214),
    .X(net417));
 sky130_fd_sc_hd__and2_0 c676 (.A(net403),
    .B(net414),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 c677 (.A(net544),
    .X(net419));
 sky130_fd_sc_hd__or4bb_1 c678 (.A(net414),
    .B(net1013),
    .C_N(net1001),
    .D_N(net207),
    .X(net420));
 sky130_fd_sc_hd__or4bb_1 c679 (.A(net405),
    .B(net404),
    .C_N(net1003),
    .D_N(net414),
    .X(net421));
 sky130_fd_sc_hd__and2_0 c680 (.A(net417),
    .B(net416),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 c681 (.A(net544),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net544),
    .X(net424));
 sky130_fd_sc_hd__buf_1 c683 (.A(net543),
    .X(net425));
 sky130_fd_sc_hd__and2_0 c684 (.A(net329),
    .B(net1031),
    .X(net426));
 sky130_fd_sc_hd__and3_1 c685 (.A(net106),
    .B(net325),
    .C(net1018),
    .X(net427));
 sky130_fd_sc_hd__and2_0 c686 (.A(net424),
    .B(net423),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 c687 (.A(net543),
    .X(net429));
 sky130_fd_sc_hd__and3_1 c688 (.A(net324),
    .B(net1069),
    .C(net969),
    .X(net430));
 sky130_fd_sc_hd__and3_1 c689 (.A(net426),
    .B(net994),
    .C(net427),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c690 (.A(net427),
    .B(net314),
    .C(net978),
    .X(net432));
 sky130_fd_sc_hd__and2_0 c691 (.A(net335),
    .B(net998),
    .X(net433));
 sky130_fd_sc_hd__and3_1 c692 (.A(net428),
    .B(net969),
    .C(net314),
    .X(net434));
 sky130_fd_sc_hd__and2_0 c693 (.A(net989),
    .B(net429),
    .X(net435));
 sky130_fd_sc_hd__and2_0 c694 (.A(net1001),
    .B(net433),
    .X(net436));
 sky130_fd_sc_hd__and3_1 c695 (.A(net322),
    .B(net409),
    .C(net433),
    .X(net437));
 sky130_fd_sc_hd__and3_1 c696 (.A(net416),
    .B(net1070),
    .C(net437),
    .X(net438));
 sky130_fd_sc_hd__or4bb_1 c697 (.A(net419),
    .B(net317),
    .C_N(net432),
    .D_N(net409),
    .X(net439));
 sky130_fd_sc_hd__and3_1 c698 (.A(net969),
    .B(net1014),
    .C(net425),
    .X(net440));
 sky130_fd_sc_hd__or4bb_2 c699 (.A(net435),
    .B(net305),
    .C_N(net427),
    .D_N(net439),
    .X(net441));
 sky130_fd_sc_hd__and3_1 c700 (.A(net1008),
    .B(net120),
    .C(net437),
    .X(net442));
 sky130_fd_sc_hd__and3_1 c701 (.A(net437),
    .B(net317),
    .C(net438),
    .X(net443));
 sky130_fd_sc_hd__and3_1 c702 (.A(net105),
    .B(net1003),
    .C(net438),
    .X(net444));
 sky130_fd_sc_hd__or4bb_1 c703 (.A(net436),
    .B(net1060),
    .C_N(net438),
    .D_N(net954),
    .X(net445));
 sky130_fd_sc_hd__and3_1 c704 (.A(net432),
    .B(net427),
    .C(net968),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net549),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 c706 (.A(net548),
    .X(net448));
 sky130_fd_sc_hd__and3_1 c707 (.A(net446),
    .B(net989),
    .C(net1007),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net613),
    .A1(net417),
    .A2(net432),
    .A3(net438),
    .S0(net310),
    .S1(net666),
    .X(net450));
 sky130_fd_sc_hd__and3_1 c709 (.A(net431),
    .B(net403),
    .C(net962),
    .X(net451));
 sky130_fd_sc_hd__and3_1 c710 (.A(net406),
    .B(net1058),
    .C(net335),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 c711 (.A(net525),
    .X(net453));
 sky130_fd_sc_hd__or4bb_1 c712 (.A(net325),
    .B(net301),
    .C_N(net1018),
    .D_N(net968),
    .X(net454));
 sky130_fd_sc_hd__and3_1 c713 (.A(net332),
    .B(net121),
    .C(net1059),
    .X(net455));
 sky130_fd_sc_hd__and3_1 c714 (.A(net422),
    .B(net425),
    .C(net1058),
    .X(net456));
 sky130_fd_sc_hd__and3_1 c715 (.A(net413),
    .B(net135),
    .C(net335),
    .X(net457));
 sky130_fd_sc_hd__and3_1 c716 (.A(net207),
    .B(net451),
    .C(net1019),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 c717 (.A(net524),
    .X(net459));
 sky130_fd_sc_hd__dlymetal6s2s_1 c718 (.A(net565),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net460),
    .A1(net430),
    .A2(net757),
    .A3(net334),
    .S0(net1016),
    .S1(net452),
    .X(net461));
 sky130_fd_sc_hd__and3_1 c720 (.A(net358),
    .B(net998),
    .C(net460),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net404),
    .A1(net448),
    .A2(net1016),
    .A3(net256),
    .S0(net990),
    .S1(net455),
    .X(net463));
 sky130_fd_sc_hd__or4bb_1 c722 (.A(net459),
    .B(net440),
    .C_N(net998),
    .D_N(net968),
    .X(net464));
 sky130_fd_sc_hd__or4bb_1 c723 (.A(net449),
    .B(net458),
    .C_N(net464),
    .D_N(net772),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net412),
    .A1(net464),
    .A2(net962),
    .A3(net1060),
    .S0(net445),
    .S1(net1022),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net315),
    .A1(net591),
    .A2(net460),
    .A3(net458),
    .S0(net532),
    .S1(net1022),
    .X(net467));
 sky130_fd_sc_hd__and3_1 c726 (.A(net1010),
    .B(net439),
    .C(net1059),
    .X(net468));
 sky130_fd_sc_hd__or4bb_1 c727 (.A(net263),
    .B(net591),
    .C_N(net1052),
    .D_N(net578),
    .X(net469));
 sky130_fd_sc_hd__a2111o_1 c728 (.A1(net305),
    .A2(net268),
    .B1(net341),
    .C1(net953),
    .D1(net355),
    .X(net470));
 sky130_fd_sc_hd__sdfrbp_1 c729 (.CLK(clknet_2_0__leaf_clk),
    .D(net415),
    .RESET_B(net367),
    .SCD(net1007),
    .SCE(net434),
    .Q(net472),
    .Q_N(net471));
 sky130_fd_sc_hd__or4bb_1 c730 (.A(net771),
    .B(net438),
    .C_N(net367),
    .D_N(net716),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net271),
    .A1(net953),
    .A2(net471),
    .A3(net1056),
    .S0(net632),
    .S1(net355),
    .X(net474));
 sky130_fd_sc_hd__or4bb_1 c732 (.A(net50),
    .B(net1036),
    .C_N(net305),
    .D_N(net972),
    .X(net475));
 sky130_fd_sc_hd__or4bb_2 c733 (.A(net345),
    .B(net442),
    .C_N(net968),
    .D_N(net1018),
    .X(net476));
 sky130_fd_sc_hd__and3_1 c734 (.A(net1007),
    .B(net1069),
    .C(net765),
    .X(net477));
 sky130_fd_sc_hd__or4bb_1 c735 (.A(net350),
    .B(net1007),
    .C_N(net535),
    .D_N(net1023),
    .X(net478));
 sky130_fd_sc_hd__or4bb_1 c736 (.A(net478),
    .B(net230),
    .C_N(net1003),
    .D_N(net549),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net472),
    .A1(net445),
    .A2(net954),
    .A3(net977),
    .S0(net462),
    .S1(net998),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net420),
    .A1(net434),
    .A2(net172),
    .A3(net1067),
    .S0(net765),
    .S1(net1022),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 c739 (.A(net566),
    .X(net482));
 sky130_fd_sc_hd__or4bb_1 c740 (.A(net172),
    .B(net1056),
    .C_N(net1006),
    .D_N(net530),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net379),
    .A1(net468),
    .A2(net1069),
    .A3(net462),
    .S0(net757),
    .S1(net476),
    .X(net484));
 sky130_fd_sc_hd__or4bb_1 c742 (.A(net370),
    .B(net453),
    .C_N(net482),
    .D_N(net977),
    .X(net485));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(net115),
    .A2(net84),
    .B1(net225),
    .C1(net574),
    .D1(net462),
    .X(net665));
 sky130_fd_sc_hd__a2111o_1 c744 (.A1(net611),
    .A2(net479),
    .B1(net84),
    .C1(net954),
    .D1(net476),
    .X(net486));
 sky130_fd_sc_hd__or4bb_1 c745 (.A(net485),
    .B(net958),
    .C_N(net554),
    .D_N(net1023),
    .X(net487));
 sky130_fd_sc_hd__or4bb_1 c746 (.A(net456),
    .B(net450),
    .C_N(net487),
    .D_N(net529),
    .X(net488));
 sky130_fd_sc_hd__sdfbbp_1 c747 (.CLK(clknet_2_3__leaf_clk),
    .D(net296),
    .RESET_B(net483),
    .SCD(net972),
    .SCE(net266),
    .SET_B(net555),
    .Q(net490),
    .Q_N(net489));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net341),
    .A1(net598),
    .A2(net386),
    .A3(net1020),
    .S0(net1016),
    .S1(net716),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net447),
    .A1(net1030),
    .A2(net363),
    .A3(net402),
    .S0(net490),
    .S1(net1051),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c750 (.A0(net108),
    .A1(net977),
    .A2(net394),
    .A3(net1070),
    .S0(net533),
    .S1(net716),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net266),
    .A1(net307),
    .A2(net596),
    .A3(net1018),
    .S0(net441),
    .S1(net553),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net470),
    .A1(net359),
    .A2(net387),
    .A3(net587),
    .S0(net568),
    .S1(net773),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net632),
    .A1(net474),
    .A2(net1052),
    .A3(net489),
    .S0(net542),
    .S1(net1023),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net1049),
    .A1(net1014),
    .A2(net477),
    .A3(net492),
    .S0(net1067),
    .S1(net1018),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net998),
    .A1(net1051),
    .A2(net964),
    .A3(net560),
    .S0(clknet_1_1__leaf_net561),
    .S1(clknet_1_0__leaf_net562),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net986),
    .A1(net641),
    .A2(net122),
    .A3(net498),
    .S0(net1032),
    .S1(clknet_1_0__leaf_net561),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net284),
    .A1(net347),
    .A2(net225),
    .A3(net380),
    .S0(net681),
    .S1(net972),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net210),
    .A1(net351),
    .A2(net392),
    .A3(net998),
    .S0(net1051),
    .S1(net558),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net491),
    .A1(net136),
    .A2(net469),
    .A3(net500),
    .S0(net355),
    .S1(clknet_1_1__leaf_net562),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net441),
    .A1(net256),
    .A2(net399),
    .A3(net398),
    .S0(net977),
    .S1(net210),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net957),
    .A1(net457),
    .A2(net499),
    .A3(net502),
    .S0(net1049),
    .S1(net535),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net411),
    .A1(net685),
    .A2(net378),
    .A3(net641),
    .S0(net1023),
    .S1(clknet_1_1__leaf_net563),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net757),
    .A1(net462),
    .A2(net475),
    .A3(net490),
    .S0(net36),
    .S1(clknet_1_0__leaf_net563),
    .X(net506));
 sky130_fd_sc_hd__mux4_2 c764 (.A0(net994),
    .A1(net391),
    .A2(net493),
    .A3(net590),
    .S0(net398),
    .S1(net545),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(clknet_1_0__leaf_net506),
    .A1(net1051),
    .A2(net1016),
    .A3(net396),
    .S0(net210),
    .S1(net574),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net279),
    .A1(net355),
    .A2(net590),
    .A3(net136),
    .S0(net681),
    .S1(net555),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(net454),
    .A1(net501),
    .A2(net509),
    .A3(net968),
    .S0(net546),
    .S1(net1023),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net505),
    .A1(net275),
    .A2(net377),
    .A3(net587),
    .S0(clknet_1_1__leaf_net506),
    .X(net511));
 sky130_fd_sc_hd__mux4_2 c769 (.A0(net342),
    .A1(net280),
    .A2(net510),
    .A3(net507),
    .S0(net545),
    .S1(net551),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net506 (.A(net506),
    .X(clknet_0_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_0__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net506 (.A(clknet_0_net506),
    .X(clknet_1_1__leaf_net506));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clone10 (.A(net761),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 clone20 (.A(net1033),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 fanout175 (.A(net968),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 fanout176 (.A(net707),
    .X(net741));
 sky130_fd_sc_hd__buf_1 fanout177 (.A(net972),
    .X(net742));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net667),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 fanout179 (.A(net119),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 fanout180 (.A(net119),
    .X(net745));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(net1033),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 fanout182 (.A(net588),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net1022),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net560),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net1024),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net539),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net400),
    .X(net776));
 sky130_fd_sc_hd__buf_2 input1 (.A(net777),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(net786),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(net787),
    .X(net576));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(net788),
    .X(net577));
 sky130_fd_sc_hd__buf_2 input13 (.A(net789),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(net790),
    .X(net579));
 sky130_fd_sc_hd__buf_1 input15 (.A(net791),
    .X(net580));
 sky130_fd_sc_hd__buf_2 input16 (.A(net792),
    .X(net581));
 sky130_fd_sc_hd__buf_1 input17 (.A(net793),
    .X(net582));
 sky130_fd_sc_hd__buf_2 input18 (.A(net794),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(net795),
    .X(net584));
 sky130_fd_sc_hd__buf_1 input2 (.A(net778),
    .X(net550));
 sky130_fd_sc_hd__buf_1 input20 (.A(net796),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(net797),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(net798),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net799),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(net800),
    .X(net589));
 sky130_fd_sc_hd__buf_1 input25 (.A(net801),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(net802),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net803),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(net804),
    .X(net593));
 sky130_fd_sc_hd__buf_1 input29 (.A(net805),
    .X(net594));
 sky130_fd_sc_hd__buf_6 input3 (.A(net779),
    .X(net568));
 sky130_fd_sc_hd__buf_2 input30 (.A(net806),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(net807),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(net808),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(net809),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(net810),
    .X(net599));
 sky130_fd_sc_hd__buf_4 input35 (.A(net811),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(net812),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(net813),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(net814),
    .X(net603));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(net815),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net780),
    .X(net569));
 sky130_fd_sc_hd__buf_1 input40 (.A(net816),
    .X(net605));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(net817),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(net818),
    .X(net607));
 sky130_fd_sc_hd__buf_1 input43 (.A(net819),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(net820),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net821),
    .X(net610));
 sky130_fd_sc_hd__buf_2 input46 (.A(net822),
    .X(net611));
 sky130_fd_sc_hd__buf_1 input47 (.A(net823),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(net824),
    .X(net613));
 sky130_fd_sc_hd__buf_1 input49 (.A(net825),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(net781),
    .X(net570));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(net826),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(net827),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net828),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(net829),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net830),
    .X(net619));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(net831),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(net832),
    .X(net621));
 sky130_fd_sc_hd__buf_1 input57 (.A(net833),
    .X(net622));
 sky130_fd_sc_hd__buf_2 input58 (.A(net834),
    .X(net623));
 sky130_fd_sc_hd__buf_1 input59 (.A(net835),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net782),
    .X(net571));
 sky130_fd_sc_hd__buf_1 input60 (.A(net836),
    .X(net625));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(net837),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(net838),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(net839),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net840),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(net841),
    .X(net630));
 sky130_fd_sc_hd__buf_1 input66 (.A(net842),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(net843),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(net844),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(net845),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(net783),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(net846),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(net847),
    .X(net636));
 sky130_fd_sc_hd__buf_1 input72 (.A(net848),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(net849),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(net850),
    .X(net639));
 sky130_fd_sc_hd__buf_1 input75 (.A(net851),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(net852),
    .X(net641));
 sky130_fd_sc_hd__buf_1 input77 (.A(net853),
    .X(net642));
 sky130_fd_sc_hd__buf_1 input78 (.A(net854),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(net855),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(net784),
    .X(net573));
 sky130_fd_sc_hd__buf_1 input80 (.A(net856),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(net857),
    .X(net646));
 sky130_fd_sc_hd__buf_1 input82 (.A(net858),
    .X(net647));
 sky130_fd_sc_hd__buf_1 input83 (.A(net859),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(net860),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(net861),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(net862),
    .X(net651));
 sky130_fd_sc_hd__buf_1 input87 (.A(net863),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net864),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(net865),
    .X(net654));
 sky130_fd_sc_hd__buf_2 input9 (.A(net785),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(net866),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(net867),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(net868),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(net869),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(net870),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(net871),
    .X(net660));
 sky130_fd_sc_hd__buf_1 input96 (.A(net872),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(net873),
    .X(net662));
 sky130_fd_sc_hd__buf_2 input98 (.A(net874),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(net875),
    .X(net664));
 sky130_fd_sc_hd__a2111o_1 merge782 (.A1(net418),
    .A2(net303),
    .B1(net421),
    .C1(net411),
    .D1(net422),
    .X(net513));
 sky130_fd_sc_hd__or4bb_1 merge783 (.A(net167),
    .B(net752),
    .C_N(net145),
    .D_N(net175),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 merge784 (.A0(net99),
    .A1(net418),
    .A2(net217),
    .A3(net406),
    .S0(net420),
    .S1(net760),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net281),
    .A1(net192),
    .A2(net189),
    .A3(net288),
    .S0(net195),
    .S1(net276),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 merge786 (.A0(net357),
    .A1(net616),
    .A2(net352),
    .A3(net164),
    .S0(net764),
    .S1(net972),
    .X(net517));
 sky130_fd_sc_hd__or4bb_1 merge787 (.A(net595),
    .B(net175),
    .C_N(net176),
    .D_N(net966),
    .X(net518));
 sky130_fd_sc_hd__a2111o_4 merge788 (.A1(net344),
    .A2(net338),
    .B1(net328),
    .C1(net216),
    .X(net540));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net407),
    .A1(net334),
    .A2(net613),
    .A3(net443),
    .S0(net954),
    .S1(net1077),
    .X(net520));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net258),
    .A1(net686),
    .A2(net641),
    .A3(net222),
    .S0(net260),
    .S1(net632),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net425),
    .A1(net407),
    .A2(net415),
    .A3(net206),
    .S0(net762),
    .S1(net1063),
    .X(net522));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net147),
    .A1(net360),
    .A2(net676),
    .A3(net591),
    .S0(net365),
    .S1(net1065),
    .X(net523));
 sky130_fd_sc_hd__sdfbbn_1 merge793 (.CLK_N(clknet_2_0__leaf_clk),
    .D(net252),
    .RESET_B(net106),
    .SCD(net587),
    .SCE(net452),
    .SET_B(net444),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net191),
    .A1(net660),
    .A2(net742),
    .A3(net180),
    .S0(net575),
    .S1(net663),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net455),
    .A1(net312),
    .A2(net951),
    .A3(net193),
    .S0(net282),
    .S1(net290),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net1005),
    .A1(net216),
    .A2(net763),
    .A3(net237),
    .S0(net476),
    .S1(net457),
    .X(net528));
 sky130_fd_sc_hd__dfrbp_1 merge797 (.CLK(clknet_2_3__leaf_clk),
    .D(net373),
    .RESET_B(net369),
    .Q(net530),
    .Q_N(net529));
 sky130_fd_sc_hd__and2_0 merge798 (.A(net197),
    .B(net526),
    .X(net531));
 sky130_fd_sc_hd__dfrbp_1 merge799 (.CLK(clknet_2_0__leaf_clk),
    .D(net461),
    .RESET_B(net465),
    .Q(net533),
    .Q_N(net532));
 sky130_fd_sc_hd__and2_0 merge800 (.A(net514),
    .B(net521),
    .X(net534));
 sky130_fd_sc_hd__dfrtn_1 merge801 (.CLK_N(clknet_2_1__leaf_clk),
    .D(net473),
    .RESET_B(net480),
    .Q(net535));
 sky130_fd_sc_hd__and2_4 merge802 (.A(net512),
    .B(net494),
    .X(net536));
 sky130_fd_sc_hd__and2_0 merge803 (.A(net515),
    .B(net522),
    .X(net537));
 sky130_fd_sc_hd__and2_0 merge804 (.A(net287),
    .B(net295),
    .X(net538));
 sky130_fd_sc_hd__dfrtp_1 merge805 (.CLK(clknet_2_2__leaf_clk),
    .D(net382),
    .RESET_B(net383),
    .Q(net539));
 sky130_fd_sc_hd__dfrtp_4 merge806 (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net337),
    .Q(net540));
 sky130_fd_sc_hd__dfrtp_1 merge807 (.CLK(clknet_2_2__leaf_clk),
    .D(net518),
    .RESET_B(net531),
    .Q(net714));
 sky130_fd_sc_hd__dfsbp_2 merge808 (.CLK(clknet_2_2__leaf_clk),
    .D(net294),
    .SET_B(net516),
    .Q(net542),
    .Q_N(net541));
 sky130_fd_sc_hd__dfsbp_1 merge809 (.CLK(clknet_2_0__leaf_clk),
    .D(net513),
    .SET_B(net537),
    .Q(net544),
    .Q_N(net543));
 sky130_fd_sc_hd__dfstp_1 merge810 (.CLK(clknet_2_3__leaf_clk),
    .D(net536),
    .SET_B(net495),
    .Q(net545));
 sky130_fd_sc_hd__dfstp_1 merge811 (.CLK(clknet_2_3__leaf_clk),
    .D(net384),
    .SET_B(net385),
    .Q(net546));
 sky130_fd_sc_hd__dfstp_2 merge812 (.CLK(clknet_2_3__leaf_clk),
    .D(net517),
    .SET_B(net523),
    .Q(net547));
 sky130_fd_sc_hd__dlrbn_1 merge813 (.D(net466),
    .GATE_N(clknet_2_0__leaf_clk),
    .RESET_B(net520),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__dlrbn_1 merge814 (.GATE_N(clknet_2_3__leaf_clk),
    .RESET_B(net508),
    .Q(net551),
    .Q_N(net511));
 sky130_fd_sc_hd__dlrbp_1 merge815 (.D(net538),
    .GATE(clknet_2_2__leaf_clk),
    .RESET_B(net534),
    .Q(net680),
    .Q_N(net552));
 sky130_fd_sc_hd__dlrbp_1 merge816 (.D(net481),
    .GATE(clknet_2_1__leaf_clk),
    .RESET_B(net486),
    .Q(net554),
    .Q_N(net553));
 sky130_fd_sc_hd__dlrtn_1 merge817 (.D(net488),
    .GATE_N(clknet_2_1__leaf_clk),
    .RESET_B(net504),
    .Q(net555));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net665),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net666),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net972),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net668),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net669),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net670),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net671),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net672),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net673),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net674),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net675),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net676),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net677),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net678),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net679),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net680),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net1003),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net992),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net683),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net684),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net1000),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net686),
    .X(net897));
 sky130_fd_sc_hd__buf_1 output122 (.A(net687),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net688),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net689),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net690),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net691),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net692),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net693),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net694),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net695),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net696),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net1026),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net956),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net1040),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net700),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net701),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net702),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net703),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net704),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net705),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net706),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net967),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net708),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net709),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net710),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net711),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net712),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net1028),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net714),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net715),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net716),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net717),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net718),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net719),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net720),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net721),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net722),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net964),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net724),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net725),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net1027),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net727),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net728),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net1021),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net730),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net731),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net1019),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net733),
    .X(net944));
 sky130_fd_sc_hd__buf_1 output169 (.A(net734),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net735),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net736),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net737),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net1038),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net739),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(net1071),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer11 (.A(net1072),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(net1082),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(net1077),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(net1082),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(net344),
    .X(net762));
 sky130_fd_sc_hd__buf_1 rebuffer16 (.A(net1081),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 rebuffer17 (.A(net763),
    .X(net764));
 sky130_fd_sc_hd__buf_1 rebuffer18 (.A(net953),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(net765),
    .X(net766));
 sky130_fd_sc_hd__buf_1 rebuffer2 (.A(net1074),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer21 (.A(net66),
    .X(net768));
 sky130_fd_sc_hd__buf_1 rebuffer22 (.A(net1073),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(net769),
    .X(net770));
 sky130_fd_sc_hd__buf_1 rebuffer24 (.A(net14),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(net749),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(net247),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net1078),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(net752),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer7 (.A(net59),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(net394),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer9 (.A(net758),
    .X(net756));
 sky130_fd_sc_hd__dfxbp_1 s818 (.CLK(clknet_2_2__leaf_clk),
    .D(net375),
    .Q(net557),
    .Q_N(net556));
 sky130_fd_sc_hd__dfxbp_1 s819 (.CLK(clknet_2_3__leaf_clk),
    .D(net401),
    .Q(net558));
 sky130_fd_sc_hd__dfxtp_1 s820 (.CLK(clknet_2_0__leaf_clk),
    .D(net463),
    .Q(net559));
 sky130_fd_sc_hd__dfxtp_2 s821 (.CLK(clknet_2_1__leaf_clk),
    .D(net467),
    .Q(net716));
 sky130_fd_sc_hd__dfxtp_1 s822 (.CLK(clknet_2_1__leaf_clk),
    .D(net484),
    .Q(net560));
 sky130_fd_sc_hd__dlclkp_1 s823 (.CLK(clknet_2_1__leaf_clk),
    .GATE(net496),
    .GCLK(net561));
 sky130_fd_sc_hd__dlclkp_2 s824 (.CLK(clknet_2_1__leaf_clk),
    .GATE(net497),
    .GCLK(net562));
 sky130_fd_sc_hd__dlclkp_4 s825 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net503),
    .GCLK(net563));
 sky130_fd_sc_hd__dlxbn_1 s826 (.D(net527),
    .GATE_N(clknet_2_0__leaf_clk),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__dlxbn_1 s827 (.D(net528),
    .GATE_N(clknet_2_1__leaf_clk),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(in0),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(in1),
    .X(net778));
 sky130_fd_sc_hd__buf_1 input102 (.A(in10),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(in11),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(in12),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(in13),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(in14),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(in15),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(in16),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(in17),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(in18),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(in19),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(in2),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(in20),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(in21),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(in22),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(in23),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(in24),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(in25),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(in26),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(in27),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(in28),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(in29),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(in3),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(in30),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(in31),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(in32),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(in33),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(in34),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(in35),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(in36),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(in37),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(in38),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(in39),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(in4),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(in40),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(in41),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(in42),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(in43),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(in44),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(in45),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(in46),
    .X(net818));
 sky130_fd_sc_hd__buf_1 input142 (.A(in47),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(in48),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(in49),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(in5),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(in50),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(in51),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(in52),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(in53),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(in54),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(in55),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(in56),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(in57),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(in58),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(in59),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(in6),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(in60),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(in61),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(in62),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(in63),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(in64),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(in65),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(in66),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(in67),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(in68),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(in69),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(in7),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(in70),
    .X(net845));
 sky130_fd_sc_hd__dlymetal6s2s_1 input169 (.A(in71),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(in72),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(in73),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(in74),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(in75),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(in76),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(in77),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(in78),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(in79),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(in8),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(in80),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(in81),
    .X(net857));
 sky130_fd_sc_hd__buf_1 input181 (.A(in82),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(in83),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(in84),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(in85),
    .X(net861));
 sky130_fd_sc_hd__buf_1 input185 (.A(in86),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(in87),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(in88),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(in89),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(in9),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(in90),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(in91),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(in92),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(in93),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(in94),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(in95),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(in97),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(in98),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(in99),
    .X(net875));
 sky130_fd_sc_hd__buf_2 output199 (.A(net876),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output200 (.A(net877),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output201 (.A(net878),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output202 (.A(net879),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output203 (.A(net880),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output204 (.A(net881),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output205 (.A(net882),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output206 (.A(net883),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output207 (.A(net884),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output208 (.A(net885),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output209 (.A(net886),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output210 (.A(net887),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output211 (.A(net888),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output212 (.A(net889),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output213 (.A(net890),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output214 (.A(net891),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output215 (.A(net892),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output216 (.A(net893),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output217 (.A(net894),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output218 (.A(net895),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output219 (.A(net896),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output220 (.A(net897),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output221 (.A(net898),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output222 (.A(net899),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output223 (.A(net900),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output224 (.A(net901),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output225 (.A(net902),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output226 (.A(net903),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_4 output227 (.A(net904),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output228 (.A(net905),
    .X(out46));
 sky130_fd_sc_hd__clkbuf_4 output229 (.A(net906),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output230 (.A(net907),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output231 (.A(net908),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_4 output232 (.A(net909),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output233 (.A(net910),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output234 (.A(net911),
    .X(out52));
 sky130_fd_sc_hd__clkbuf_4 output235 (.A(net912),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output236 (.A(net913),
    .X(out54));
 sky130_fd_sc_hd__clkbuf_4 output237 (.A(net914),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output238 (.A(net915),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output239 (.A(net916),
    .X(out58));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net917),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output241 (.A(net918),
    .X(out6));
 sky130_fd_sc_hd__clkbuf_4 output242 (.A(net919),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output243 (.A(net920),
    .X(out61));
 sky130_fd_sc_hd__clkbuf_4 output244 (.A(net921),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_4 output245 (.A(net922),
    .X(out63));
 sky130_fd_sc_hd__clkbuf_4 output246 (.A(net923),
    .X(out65));
 sky130_fd_sc_hd__buf_2 output247 (.A(net924),
    .X(out67));
 sky130_fd_sc_hd__clkbuf_4 output248 (.A(net925),
    .X(out68));
 sky130_fd_sc_hd__clkbuf_4 output249 (.A(net926),
    .X(out69));
 sky130_fd_sc_hd__buf_2 output250 (.A(net927),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output251 (.A(net928),
    .X(out71));
 sky130_fd_sc_hd__clkbuf_4 output252 (.A(net929),
    .X(out72));
 sky130_fd_sc_hd__buf_2 output253 (.A(net930),
    .X(out73));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net931),
    .X(out75));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net932),
    .X(out76));
 sky130_fd_sc_hd__clkbuf_4 output256 (.A(net933),
    .X(out79));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net934),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output258 (.A(net935),
    .X(out81));
 sky130_fd_sc_hd__buf_2 output259 (.A(net936),
    .X(out82));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net937),
    .X(out83));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net938),
    .X(out84));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net939),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output263 (.A(net940),
    .X(out86));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net941),
    .X(out88));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net942),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output266 (.A(net943),
    .X(out9));
 sky130_fd_sc_hd__buf_2 output267 (.A(net944),
    .X(out91));
 sky130_fd_sc_hd__buf_2 output268 (.A(net945),
    .X(out92));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net946),
    .X(out93));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net947),
    .X(out94));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net948),
    .X(out95));
 sky130_fd_sc_hd__buf_2 output272 (.A(net949),
    .X(out96));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net950),
    .X(out98));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout274 (.A(net349),
    .X(net951));
 sky130_fd_sc_hd__buf_6 fanout275 (.A(net540),
    .X(net952));
 sky130_fd_sc_hd__buf_6 fanout276 (.A(net255),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net442),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net698),
    .X(net955));
 sky130_fd_sc_hd__buf_1 fanout279 (.A(net698),
    .X(net956));
 sky130_fd_sc_hd__buf_2 fanout280 (.A(net188),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net76),
    .X(net958));
 sky130_fd_sc_hd__buf_1 fanout282 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout283 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(net740),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_2 fanout285 (.A(net307),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 fanout286 (.A(net233),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net723),
    .X(net964));
 sky130_fd_sc_hd__buf_1 fanout288 (.A(net742),
    .X(net965));
 sky130_fd_sc_hd__buf_2 fanout289 (.A(net742),
    .X(net966));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout291 (.A(net741),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_2 fanout292 (.A(net227),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(net226),
    .X(net970));
 sky130_fd_sc_hd__buf_1 fanout294 (.A(net743),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(net743),
    .X(net972));
 sky130_fd_sc_hd__buf_1 fanout296 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_1 fanout297 (.A(net221),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_2 fanout298 (.A(net155),
    .X(net975));
 sky130_fd_sc_hd__buf_1 fanout299 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_2 fanout300 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_2 fanout301 (.A(net745),
    .X(net978));
 sky130_fd_sc_hd__buf_1 fanout302 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_2 fanout304 (.A(net744),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(net147),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_2 fanout306 (.A(net201),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(net129),
    .X(net984));
 sky130_fd_sc_hd__buf_2 fanout308 (.A(net116),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_2 fanout309 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net112),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(net126),
    .X(net988));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout312 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(net110),
    .X(net990));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout314 (.A(net711),
    .X(net991));
 sky130_fd_sc_hd__buf_2 fanout315 (.A(net682),
    .X(net992));
 sky130_fd_sc_hd__buf_6 fanout316 (.A(net43),
    .X(net993));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(net28),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net132),
    .X(net995));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout319 (.A(net57),
    .X(net996));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout320 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(net44),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(net29),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_2 fanout323 (.A(net685),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(net300),
    .X(net1001));
 sky130_fd_sc_hd__buf_1 fanout325 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout326 (.A(net681),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_2 fanout327 (.A(net120),
    .X(net1004));
 sky130_fd_sc_hd__buf_2 fanout328 (.A(net42),
    .X(net1005));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(net40),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 fanout330 (.A(net40),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 fanout331 (.A(net36),
    .X(net1008));
 sky130_fd_sc_hd__buf_1 fanout332 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(net23),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_2 fanout334 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout335 (.A(net21),
    .X(net1012));
 sky130_fd_sc_hd__buf_1 fanout336 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__buf_2 fanout337 (.A(net20),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(net108),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(net60),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 fanout340 (.A(net34),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_2 fanout341 (.A(net34),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 fanout342 (.A(net732),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net732),
    .X(net1020));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout344 (.A(net729),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__buf_2 fanout346 (.A(net559),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_2 fanout347 (.A(net714),
    .X(net1024));
 sky130_fd_sc_hd__buf_8 fanout348 (.A(net746),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(net697),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net726),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout351 (.A(net713),
    .X(net1028));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout352 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_4 fanout353 (.A(net19),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(net17),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net17),
    .X(net1032));
 sky130_fd_sc_hd__buf_8 fanout356 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__buf_6 fanout357 (.A(net747),
    .X(net1034));
 sky130_fd_sc_hd__buf_1 fanout358 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(net104),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_2 fanout360 (.A(net15),
    .X(net1037));
 sky130_fd_sc_hd__buf_1 fanout361 (.A(net738),
    .X(net1038));
 sky130_fd_sc_hd__buf_1 fanout362 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(net699),
    .X(net1040));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout364 (.A(net660),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(net655),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(net574),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_2 fanout367 (.A(net573),
    .X(net1044));
 sky130_fd_sc_hd__buf_2 fanout368 (.A(net644),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_2 fanout369 (.A(net572),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 fanout370 (.A(net571),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_2 fanout371 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_4 fanout372 (.A(net622),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_4 fanout374 (.A(net617),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net612),
    .X(net1052));
 sky130_fd_sc_hd__buf_1 fanout376 (.A(net612),
    .X(net1053));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net611),
    .X(net1054));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout378 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net569),
    .X(net1056));
 sky130_fd_sc_hd__buf_6 fanout380 (.A(net600),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_4 fanout381 (.A(net598),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net596),
    .X(net1059));
 sky130_fd_sc_hd__buf_6 fanout383 (.A(net568),
    .X(net1060));
 sky130_fd_sc_hd__buf_2 fanout384 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net592),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net589),
    .X(net1063));
 sky130_fd_sc_hd__buf_1 fanout387 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__buf_4 fanout388 (.A(net585),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net550),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout391 (.A(net580),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_2 fanout392 (.A(net578),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(net576),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net63),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net32),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net45),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net59),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1074),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net255),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net952),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net247),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net1034),
    .X(net1079));
 sky130_fd_sc_hd__buf_2 rebuffer32 (.A(net1079),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net344),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net540),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net255),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net43),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net1034),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net746),
    .X(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0_1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X_1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_B_1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_X_1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B_1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A_1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_B_1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X_1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_C_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0_1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X_1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X_1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1_1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X_1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_C_1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B_1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_C_1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_X_1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B_1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0_1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A_1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X_1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_C_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_D (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B_1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X_1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0_1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X_1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_C_N (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_C (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_X (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X_1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone36_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B_1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X_1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_C (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_Q_1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_X_1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0_1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X_1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_C_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_RESET_B_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X_1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A_1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A_1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A_1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X_1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S0_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_C1_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S1_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X_1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_B_1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X_1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A_1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B_1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_D_N_1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X_1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0_1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X_1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A2 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2_1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X_1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1_1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X_1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_C_1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A_1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A_1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X_1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_B_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X_1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_C_1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X_1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_X (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X_1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_X (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_B (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_Q (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_B (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S0_1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0_1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X_1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_C_1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B_1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_D1_1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X_1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_C_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X_1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_X (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_X (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S0 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A1_1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X_1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_C_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_C_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X_1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_X (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X_1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_X (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_X (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_B (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone20_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_C (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_C_N (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer22_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_C (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_C1_1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A_1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A_1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1_1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B_1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_B1_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_D_N_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_D1_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_C_1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_S1_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_SCD_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_D_N_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_D_N_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_RESET_B_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A_1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_D_N_1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D_N_1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_C1_1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_C_1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_C_1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_C_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_D_N_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_D1_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_C1_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3_1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2_1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1_1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B_1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C_1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0_1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1_1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B_1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B_1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A_1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_C_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A0_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_C_N_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_D_N_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S1_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3_1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B_1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A_1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B_1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_C_N_1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3_1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_C_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_C1_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A0_1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_C_1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0_1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3_1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2_1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A_1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_B_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_C_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_C_N_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A_1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_S1_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_C_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_D1_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1_1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_SCD_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_C_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_C_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0_1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_B1_1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_B_1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3_1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0_1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B_1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_X (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_D1_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_C_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_C_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1_1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3_1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1_1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3_1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0_1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B_1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A_1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A_1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer34_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net994));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_622 ();
endmodule
