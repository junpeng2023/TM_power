module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net886;
 wire clknet_1_0__leaf_net886;
 wire clknet_1_1__leaf_net886;
 wire clknet_0_net885;
 wire clknet_1_0__leaf_net885;
 wire clknet_1_1__leaf_net885;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net961;
 wire clknet_1_0__leaf_net961;
 wire clknet_1_1__leaf_net961;
 wire clknet_0_net477;
 wire clknet_1_0__leaf_net477;
 wire clknet_1_1__leaf_net477;
 wire clknet_0_net579;
 wire clknet_1_0__leaf_net579;
 wire clknet_1_1__leaf_net579;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net476;
 wire clknet_1_0__leaf_net476;
 wire clknet_1_1__leaf_net476;
 wire clknet_0_net491;
 wire clknet_1_0__leaf_net491;
 wire clknet_1_1__leaf_net491;
 wire clknet_0_net867;
 wire clknet_1_0__leaf_net867;
 wire clknet_1_1__leaf_net867;
 wire clknet_0_net500;
 wire clknet_1_0__leaf_net500;
 wire clknet_1_1__leaf_net500;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net866;
 wire clknet_1_0__leaf_net866;
 wire clknet_1_1__leaf_net866;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net847;
 wire clknet_1_0__leaf_net847;
 wire clknet_1_1__leaf_net847;
 wire clknet_0_net358;
 wire clknet_1_0__leaf_net358;
 wire clknet_1_1__leaf_net358;
 wire clknet_0_net792;
 wire clknet_1_0__leaf_net792;
 wire clknet_1_1__leaf_net792;
 wire clknet_0_net355;
 wire clknet_1_0__leaf_net355;
 wire clknet_1_1__leaf_net355;
 wire clknet_0_net350;
 wire clknet_1_0__leaf_net350;
 wire clknet_1_1__leaf_net350;
 wire clknet_0_net353;
 wire clknet_1_0__leaf_net353;
 wire clknet_1_1__leaf_net353;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net354;
 wire clknet_1_0__leaf_net354;
 wire clknet_1_1__leaf_net354;
 wire clknet_0_net846;
 wire clknet_1_0__leaf_net846;
 wire clknet_1_1__leaf_net846;
 wire clknet_0_net588;
 wire clknet_1_0__leaf_net588;
 wire clknet_1_1__leaf_net588;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net845;
 wire clknet_1_0__leaf_net845;
 wire clknet_1_1__leaf_net845;
 wire clknet_0_net451;
 wire clknet_1_0__leaf_net451;
 wire clknet_1_1__leaf_net451;
 wire clknet_0_net455;
 wire clknet_1_0__leaf_net455;
 wire clknet_1_1__leaf_net455;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net828;
 wire clknet_1_0__leaf_net828;
 wire clknet_1_1__leaf_net828;
 wire clknet_0_net223;
 wire clknet_1_0__leaf_net223;
 wire clknet_1_1__leaf_net223;
 wire clknet_0_net254;
 wire clknet_1_0__leaf_net254;
 wire clknet_1_1__leaf_net254;
 wire clknet_0_net228;
 wire clknet_1_0__leaf_net228;
 wire clknet_1_1__leaf_net228;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net225;
 wire clknet_1_0__leaf_net225;
 wire clknet_1_1__leaf_net225;
 wire clknet_0_net748;
 wire clknet_1_0__leaf_net748;
 wire clknet_1_1__leaf_net748;
 wire clknet_0_net130;
 wire clknet_1_0__leaf_net130;
 wire clknet_1_1__leaf_net130;
 wire clknet_0_net125;
 wire clknet_1_0__leaf_net125;
 wire clknet_1_1__leaf_net125;
 wire clknet_0_net271;
 wire clknet_1_0__leaf_net271;
 wire clknet_1_1__leaf_net271;
 wire clknet_0_net243;
 wire clknet_1_0__leaf_net243;
 wire clknet_1_1__leaf_net243;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net118;
 wire clknet_1_0__leaf_net118;
 wire clknet_1_1__leaf_net118;
 wire clknet_0_net131;
 wire clknet_1_0__leaf_net131;
 wire clknet_1_1__leaf_net131;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net127;
 wire clknet_1_0__leaf_net127;
 wire clknet_1_1__leaf_net127;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net119;
 wire clknet_1_0__leaf_net119;
 wire clknet_1_1__leaf_net119;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net143;
 wire clknet_1_0__leaf_net143;
 wire clknet_1_1__leaf_net143;
 wire clknet_0_net984;
 wire clknet_1_0__leaf_net984;
 wire clknet_1_1__leaf_net984;
 wire clknet_0_net404;
 wire clknet_1_0__leaf_net404;
 wire clknet_1_1__leaf_net404;
 wire clknet_0_net793;
 wire clknet_1_0__leaf_net793;
 wire clknet_1_1__leaf_net793;
 wire clknet_0_net971;
 wire clknet_1_0__leaf_net971;
 wire clknet_1_1__leaf_net971;
 wire clknet_0_net389;
 wire clknet_1_0__leaf_net389;
 wire clknet_1_1__leaf_net389;
 wire clknet_0_net381;
 wire clknet_1_0__leaf_net381;
 wire clknet_1_1__leaf_net381;
 wire clknet_0_net379;
 wire clknet_1_0__leaf_net379;
 wire clknet_1_1__leaf_net379;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net407;
 wire clknet_1_0__leaf_net407;
 wire clknet_1_1__leaf_net407;
 wire clknet_0_net966;
 wire clknet_1_0__leaf_net966;
 wire clknet_1_1__leaf_net966;
 wire clknet_0_net1006;
 wire clknet_1_0__leaf_net1006;
 wire clknet_1_1__leaf_net1006;
 wire clknet_0_net995;
 wire clknet_1_0__leaf_net995;
 wire clknet_1_1__leaf_net995;
 wire clknet_0_net965;
 wire clknet_1_0__leaf_net965;
 wire clknet_1_1__leaf_net965;
 wire clknet_0_net991;
 wire clknet_1_0__leaf_net991;
 wire clknet_1_1__leaf_net991;
 wire clknet_0_net1001;
 wire clknet_1_0__leaf_net1001;
 wire clknet_1_1__leaf_net1001;
 wire clknet_0_net973;
 wire clknet_1_0__leaf_net973;
 wire clknet_1_1__leaf_net973;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net164;
 wire clknet_1_0__leaf_net164;
 wire clknet_1_1__leaf_net164;
 wire clknet_0_net750;
 wire clknet_1_0__leaf_net750;
 wire clknet_1_1__leaf_net750;
 wire clknet_0_net51;
 wire clknet_1_0__leaf_net51;
 wire clknet_1_1__leaf_net51;
 wire clknet_0_net47;
 wire clknet_1_0__leaf_net47;
 wire clknet_1_1__leaf_net47;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net749;
 wire clknet_1_0__leaf_net749;
 wire clknet_1_1__leaf_net749;
 wire clknet_0_net662;
 wire clknet_1_0__leaf_net662;
 wire clknet_1_1__leaf_net662;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;

 sky130_fd_sc_hd__a21bo_1 c100 (.A1(net3),
    .A2(net28),
    .B1_N(net825),
    .X(net38));
 sky130_fd_sc_hd__sdfrbp_2 c101 (.CLK(clknet_4_4_0_clk),
    .D(net26),
    .RESET_B(net37),
    .SCD(net28),
    .SCE(net8),
    .Q(net40),
    .Q_N(net39));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net32),
    .A1(net6),
    .A2(net29),
    .A3(net40),
    .S0(net915),
    .S1(net28),
    .X(net41));
 sky130_fd_sc_hd__a21bo_1 c103 (.A1(net37),
    .A2(net29),
    .B1_N(net40),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 c104 (.A(net714),
    .X(net43));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net7),
    .A2(net30),
    .B1_N(net31),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 c106 (.A(net777),
    .X(net45));
 sky130_fd_sc_hd__buf_1 c107 (.A(net713),
    .X(net46));
 sky130_fd_sc_hd__buf_1 c108 (.A(clknet_1_0__leaf_net750),
    .X(net47));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net46),
    .A1(net44),
    .A2(clknet_1_0__leaf_net47),
    .A3(net955),
    .S0(net25),
    .S1(net997),
    .X(net48));
 sky130_fd_sc_hd__xnor2_4 c110 (.A(net37),
    .B(net1062),
    .Y(net1002));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net902),
    .B(net825),
    .Y(net1000));
 sky130_fd_sc_hd__xnor2_1 c112 (.A(net8),
    .B(net822),
    .Y(net49));
 sky130_fd_sc_hd__buf_1 c113 (.A(net701),
    .X(net50));
 sky130_fd_sc_hd__buf_1 c114 (.A(clknet_1_0__leaf_net750),
    .X(net51));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net938),
    .B(net50),
    .Y(net52));
 sky130_fd_sc_hd__xnor2_4 c116 (.A(net43),
    .B(net25),
    .Y(net53));
 sky130_fd_sc_hd__xnor2_4 c117 (.A(net0),
    .B(net53),
    .Y(net978));
 sky130_fd_sc_hd__sdfbbn_1 c118 (.CLK_N(clknet_4_5_0_clk),
    .D(clknet_1_1__leaf_net51),
    .RESET_B(net949),
    .SCD(net978),
    .SCE(net43),
    .SET_B(net825),
    .Q(net998),
    .Q_N(net54));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net50),
    .B(net1021),
    .Y(net55));
 sky130_fd_sc_hd__xnor2_1 c120 (.A(net49),
    .B(net53),
    .Y(net56));
 sky130_fd_sc_hd__xnor2_1 c121 (.A(net46),
    .B(net49),
    .Y(net988));
 sky130_fd_sc_hd__clkbuf_2 c122 (.A(net701),
    .X(net981));
 sky130_fd_sc_hd__a31o_1 c123 (.A1(net34),
    .A2(net1000),
    .A3(net50),
    .B1(net25),
    .X(net57));
 sky130_fd_sc_hd__sdfbbp_1 c124 (.CLK(clknet_4_5_0_clk),
    .D(net57),
    .RESET_B(net981),
    .SCD(net52),
    .SCE(net55),
    .SET_B(net1060),
    .Q(net1005),
    .Q_N(net58));
 sky130_fd_sc_hd__buf_1 c125 (.A(net713),
    .X(net59));
 sky130_fd_sc_hd__sdfbbn_1 c126 (.CLK_N(clknet_4_5_0_clk),
    .D(net981),
    .RESET_B(net1005),
    .SCD(net57),
    .SCE(net54),
    .SET_B(net827),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__sdfbbn_1 c127 (.CLK_N(clknet_4_5_0_clk),
    .D(net55),
    .RESET_B(net988),
    .SCD(net57),
    .SCE(net58),
    .SET_B(net1079),
    .Q(net63),
    .Q_N(net62));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net944),
    .A2(net57),
    .A3(net62),
    .A4(net981),
    .B1(clknet_1_0__leaf_net51),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c129 (.A0(net59),
    .A1(net57),
    .A2(net55),
    .A3(net58),
    .S0(net62),
    .S1(net823),
    .X(net65));
 sky130_fd_sc_hd__a41o_1 c130 (.A1(net59),
    .A2(net37),
    .A3(net28),
    .A4(net702),
    .B1(clknet_1_0__leaf_net1006),
    .X(net965));
 sky130_fd_sc_hd__sdfbbp_1 c131 (.CLK(clknet_4_5_0_clk),
    .D(net63),
    .RESET_B(net981),
    .SCD(clknet_1_1__leaf_net965),
    .SCE(net1083),
    .SET_B(clknet_1_1__leaf_net1006),
    .Q(net67),
    .Q_N(net66));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net910),
    .B(net930),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net898),
    .B(net903),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net68),
    .B(net900),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net906),
    .B(net896),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net903),
    .B(net71),
    .Y(net72));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net70),
    .B(net900),
    .Y(net73));
 sky130_fd_sc_hd__a31o_2 c138 (.A1(net71),
    .A2(net72),
    .A3(net910),
    .B1(net919),
    .X(net74));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net69),
    .B(net909),
    .Y(net75));
 sky130_fd_sc_hd__clkbuf_8 c140 (.A(net734),
    .X(net76));
 sky130_fd_sc_hd__sdfrbp_1 c141 (.CLK(clknet_4_0_0_clk),
    .D(net72),
    .RESET_B(net73),
    .SCD(net75),
    .SCE(net74),
    .Q(net78),
    .Q_N(net77));
 sky130_fd_sc_hd__xnor2_2 c142 (.A(net897),
    .B(net76),
    .Y(net79));
 sky130_fd_sc_hd__buf_1 c143 (.A(net734),
    .X(net80));
 sky130_fd_sc_hd__sdfbbn_1 c144 (.CLK_N(clknet_4_0_0_clk),
    .D(net74),
    .RESET_B(net902),
    .SCD(net80),
    .SCE(net75),
    .SET_B(net78),
    .Q(net82),
    .Q_N(net81));
 sky130_fd_sc_hd__a41o_1 c145 (.A1(net80),
    .A2(net930),
    .A3(net70),
    .A4(net81),
    .B1(net68),
    .X(net83));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net900),
    .A2(net75),
    .A3(net903),
    .A4(net899),
    .B1(net930),
    .X(net84));
 sky130_fd_sc_hd__sdfbbn_2 c147 (.CLK_N(clknet_4_0_0_clk),
    .D(net84),
    .RESET_B(net83),
    .SCD(net76),
    .SCE(net73),
    .SET_B(net1077),
    .Q(net86),
    .Q_N(net85));
 sky130_fd_sc_hd__buf_1 c148 (.A(net742),
    .X(net87));
 sky130_fd_sc_hd__a41o_1 c149 (.A1(net80),
    .A2(net86),
    .A3(net69),
    .A4(net76),
    .B1(net1038),
    .X(net88));
 sky130_fd_sc_hd__a41o_4 c150 (.A1(net905),
    .A2(net79),
    .A3(net1038),
    .A4(net88),
    .B1(net75),
    .X(net89));
 sky130_fd_sc_hd__a21bo_2 c151 (.A1(net1038),
    .A2(net88),
    .B1_N(net909),
    .X(net90));
 sky130_fd_sc_hd__sdfbbp_1 c152 (.CLK(clknet_4_0_0_clk),
    .D(net86),
    .RESET_B(net79),
    .SCD(net71),
    .SCE(net84),
    .SET_B(net1038),
    .Q(net92),
    .Q_N(net91));
 sky130_fd_sc_hd__a41o_1 c153 (.A1(net902),
    .A2(net90),
    .A3(net89),
    .A4(net88),
    .B1(net74),
    .X(net93));
 sky130_fd_sc_hd__xnor2_1 c154 (.A(net82),
    .B(net915),
    .Y(net94));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net913),
    .B(net85),
    .Y(net95));
 sky130_fd_sc_hd__a31o_2 c156 (.A1(net912),
    .A2(net95),
    .A3(net927),
    .B1(net925),
    .X(net96));
 sky130_fd_sc_hd__xnor2_1 c157 (.A(net932),
    .B(net95),
    .Y(net97));
 sky130_fd_sc_hd__clkbuf_1 c158 (.A(net743),
    .X(net98));
 sky130_fd_sc_hd__a21bo_1 c159 (.A1(net920),
    .A2(net914),
    .B1_N(net1035),
    .X(net99));
 sky130_fd_sc_hd__a31o_2 c160 (.A1(net68),
    .A2(net70),
    .A3(net1035),
    .B1(net95),
    .X(net100));
 sky130_fd_sc_hd__xnor2_1 c161 (.A(net95),
    .B(net82),
    .Y(net101));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net928),
    .A1(net83),
    .A2(net96),
    .A3(net100),
    .S0(net69),
    .S1(net1035),
    .X(net102));
 sky130_fd_sc_hd__a21bo_2 c163 (.A1(net922),
    .A2(net1035),
    .B1_N(net807),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 c164 (.A(net1063),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 c165 (.A(net709),
    .X(net105));
 sky130_fd_sc_hd__mux4_2 c166 (.A0(net925),
    .A1(net82),
    .A2(net918),
    .A3(net907),
    .S0(net91),
    .S1(net1036),
    .X(net106));
 sky130_fd_sc_hd__a21bo_1 c167 (.A1(net106),
    .A2(net96),
    .B1_N(net1035),
    .X(net107));
 sky130_fd_sc_hd__a41o_1 c168 (.A1(net105),
    .A2(net106),
    .A3(net103),
    .A4(net915),
    .B1(net1035),
    .X(net108));
 sky130_fd_sc_hd__a21bo_1 c169 (.A1(net95),
    .A2(net108),
    .B1_N(net1035),
    .X(net109));
 sky130_fd_sc_hd__sdfrtn_1 c170 (.CLK_N(clknet_4_0_0_clk),
    .D(net109),
    .RESET_B(net107),
    .SCD(net108),
    .SCE(net73),
    .Q(net110));
 sky130_fd_sc_hd__mux4_1 c171 (.A0(net108),
    .A1(net110),
    .A2(net95),
    .A3(net99),
    .S0(net106),
    .S1(net109),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net926),
    .A1(net107),
    .A2(net918),
    .A3(net108),
    .S0(net807),
    .S1(clknet_1_0__leaf_net828),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net94),
    .A1(net106),
    .A2(net99),
    .A3(net73),
    .S0(net1035),
    .S1(clknet_1_0__leaf_net828),
    .X(net113));
 sky130_fd_sc_hd__a21bo_1 c174 (.A1(net929),
    .A2(net108),
    .B1_N(clknet_1_0__leaf_net828),
    .X(net966));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net107),
    .A1(net106),
    .A2(net110),
    .A3(net1035),
    .S0(clknet_1_0__leaf_net748),
    .S1(clknet_1_0__leaf_net828),
    .X(net114));
 sky130_fd_sc_hd__xnor2_1 c176 (.A(net908),
    .B(net734),
    .Y(net115));
 sky130_fd_sc_hd__xnor2_2 c177 (.A(net939),
    .B(net942),
    .Y(net116));
 sky130_fd_sc_hd__a31o_1 c178 (.A1(net934),
    .A2(net115),
    .A3(net953),
    .B1(net733),
    .X(net117));
 sky130_fd_sc_hd__buf_1 c179 (.A(clknet_1_0__leaf_net748),
    .X(net118));
 sky130_fd_sc_hd__xnor2_1 c180 (.A(net115),
    .B(clknet_1_0__leaf_net118),
    .Y(net119));
 sky130_fd_sc_hd__sdfrtp_2 c181 (.CLK(clknet_4_1_0_clk),
    .D(net83),
    .RESET_B(net953),
    .SCD(net923),
    .SCE(net918),
    .Q(net120));
 sky130_fd_sc_hd__a31o_1 c182 (.A1(net79),
    .A2(net947),
    .A3(net100),
    .B1(net1059),
    .X(net121));
 sky130_fd_sc_hd__xnor2_2 c183 (.A(net116),
    .B(net934),
    .Y(net122));
 sky130_fd_sc_hd__a31o_2 c184 (.A1(net97),
    .A2(net948),
    .A3(net116),
    .B1(net120),
    .X(net123));
 sky130_fd_sc_hd__a21bo_1 c185 (.A1(net117),
    .A2(net1059),
    .B1_N(net69),
    .X(net124));
 sky130_fd_sc_hd__buf_1 c186 (.A(clknet_1_1__leaf_net748),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(net124),
    .A1(net1045),
    .A2(net122),
    .A3(net939),
    .S0(net1059),
    .S1(net949),
    .X(net126));
 sky130_fd_sc_hd__xnor2_1 c188 (.A(net69),
    .B(clknet_1_0__leaf_net118),
    .Y(net127));
 sky130_fd_sc_hd__xnor2_1 c189 (.A(net1),
    .B(net704),
    .Y(net128));
 sky130_fd_sc_hd__xnor2_1 c190 (.A(net128),
    .B(clknet_1_0__leaf_net118),
    .Y(net129));
 sky130_fd_sc_hd__xnor2_1 c191 (.A(clknet_1_0__leaf_net127),
    .B(clknet_1_1__leaf_net748),
    .Y(net130));
 sky130_fd_sc_hd__xnor2_1 c192 (.A(clknet_1_1__leaf_net118),
    .B(net122),
    .Y(net131));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net948),
    .A1(net122),
    .A2(clknet_1_0__leaf_net131),
    .A3(net942),
    .S0(clknet_1_0__leaf_net125),
    .S1(net128),
    .X(net132));
 sky130_fd_sc_hd__a31o_1 c194 (.A1(clknet_1_0__leaf_net131),
    .A2(net124),
    .A3(clknet_1_0__leaf_net129),
    .B1(clknet_1_0__leaf_net130),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net909),
    .A1(clknet_1_0__leaf_net129),
    .A2(net99),
    .A3(clknet_1_1__leaf_net118),
    .S0(net704),
    .S1(net829),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 c196 (.A(net963),
    .X(net135));
 sky130_fd_sc_hd__a31o_1 c197 (.A1(clknet_1_1__leaf_net130),
    .A2(net122),
    .A3(net135),
    .B1(net100),
    .X(net136));
 sky130_fd_sc_hd__buf_1 c198 (.A(net763),
    .X(net137));
 sky130_fd_sc_hd__buf_1 c199 (.A(net763),
    .X(net138));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net88),
    .A2(net103),
    .B1_N(net820),
    .X(net139));
 sky130_fd_sc_hd__a21bo_1 c201 (.A1(net137),
    .A2(clknet_1_0__leaf_net125),
    .B1_N(net1045),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 c202 (.A(net741),
    .X(net141));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net138),
    .A2(clknet_1_0__leaf_net127),
    .B1_N(clknet_1_0__leaf_net140),
    .X(net142));
 sky130_fd_sc_hd__a21bo_1 c204 (.A1(net1021),
    .A2(clknet_1_0__leaf_net119),
    .B1_N(net705),
    .X(net143));
 sky130_fd_sc_hd__dlymetal6s2s_1 c205 (.A(net763),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 c206 (.A(net763),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 c207 (.A(net747),
    .X(net146));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(net146),
    .A2(net138),
    .B1_N(clknet_1_1__leaf_net140),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net122),
    .A1(clknet_1_0__leaf_net147),
    .A2(net12),
    .A3(clknet_1_0__leaf_net125),
    .S0(net138),
    .S1(net6),
    .X(net148));
 sky130_fd_sc_hd__a31o_1 c210 (.A1(clknet_1_1__leaf_net142),
    .A2(clknet_1_1__leaf_net147),
    .A3(clknet_1_0__leaf_net143),
    .B1(net830),
    .X(net149));
 sky130_fd_sc_hd__buf_2 c211 (.A(net783),
    .X(net150));
 sky130_fd_sc_hd__a31o_2 c212 (.A1(net141),
    .A2(net103),
    .A3(net942),
    .B1(net778),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net923),
    .A1(net135),
    .A2(net151),
    .A3(net84),
    .S0(net122),
    .S1(net90),
    .X(net152));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(clknet_1_1__leaf_net127),
    .A2(net150),
    .A3(net826),
    .A4(net834),
    .B1(net835),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c215 (.A0(clknet_1_1__leaf_net153),
    .A1(net144),
    .A2(net15),
    .A3(net139),
    .S0(net923),
    .S1(net811),
    .X(net154));
 sky130_fd_sc_hd__a31o_2 c216 (.A1(net949),
    .A2(net15),
    .A3(net778),
    .B1(net835),
    .X(net155));
 sky130_fd_sc_hd__a41o_1 c217 (.A1(net12),
    .A2(clknet_1_0__leaf_net147),
    .A3(net103),
    .A4(net138),
    .B1(net835),
    .X(net156));
 sky130_fd_sc_hd__a41o_1 c218 (.A1(net155),
    .A2(clknet_1_0__leaf_net153),
    .A3(net139),
    .A4(net150),
    .B1(clknet_1_0__leaf_net143),
    .X(net157));
 sky130_fd_sc_hd__a21bo_4 c219 (.A1(net150),
    .A2(net807),
    .B1_N(net835),
    .X(net1004));
 sky130_fd_sc_hd__xnor2_1 c220 (.A(net1043),
    .B(clknet_1_1__leaf_net991),
    .Y(net158));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(clknet_1_1__leaf_net47),
    .B(net954),
    .Y(net159));
 sky130_fd_sc_hd__dlymetal6s2s_1 c222 (.A(net769),
    .X(net1009));
 sky130_fd_sc_hd__xnor2_1 c223 (.A(net957),
    .B(clknet_1_0__leaf_net47),
    .Y(net160));
 sky130_fd_sc_hd__clkbuf_1 c224 (.A(net769),
    .X(net161));
 sky130_fd_sc_hd__xnor2_1 c225 (.A(net72),
    .B(net1004),
    .Y(net162));
 sky130_fd_sc_hd__xnor2_4 c226 (.A(net1044),
    .B(net1004),
    .Y(net163));
 sky130_fd_sc_hd__a21bo_1 c227 (.A1(clknet_1_1__leaf_net158),
    .A2(net914),
    .B1_N(net163),
    .X(net164));
 sky130_fd_sc_hd__xnor2_1 c228 (.A(net163),
    .B(clknet_1_1__leaf_net147),
    .Y(net165));
 sky130_fd_sc_hd__xnor2_1 c229 (.A(clknet_1_0__leaf_net159),
    .B(clknet_1_1__leaf_net47),
    .Y(net166));
 sky130_fd_sc_hd__xnor2_4 c230 (.A(net40),
    .B(net1034),
    .Y(net167));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net954),
    .A2(net163),
    .B1_N(net167),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c232 (.A0(net167),
    .A1(net144),
    .A2(clknet_1_1__leaf_net125),
    .A3(net1034),
    .S0(net163),
    .S1(clknet_1_0__leaf_net164),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net168),
    .A1(clknet_1_0__leaf_net164),
    .A2(clknet_1_1__leaf_net159),
    .A3(net28),
    .S0(net38),
    .S1(net1034),
    .X(net170));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net38),
    .A2(net163),
    .B1_N(net167),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 c235 (.A(net741),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(net103),
    .A1(net954),
    .A2(net1013),
    .A3(net168),
    .S0(net163),
    .S1(clknet_1_0__leaf_net158),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 c237 (.A(net741),
    .X(net174));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net145),
    .A2(net710),
    .B1_N(net769),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net172),
    .A1(clknet_1_0__leaf_net165),
    .A2(net174),
    .A3(net168),
    .S0(net710),
    .S1(clknet_1_0__leaf_net991),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 c240 (.A(net760),
    .X(net177));
 sky130_fd_sc_hd__sdfbbn_1 c241 (.CLK_N(clknet_4_7_0_clk),
    .D(net177),
    .RESET_B(net168),
    .SCD(clknet_1_0__leaf_net164),
    .SCE(net834),
    .SET_B(net1073),
    .Q(net179),
    .Q_N(net178));
 sky130_fd_sc_hd__clkbuf_1 c242 (.A(net746),
    .X(net985));
 sky130_fd_sc_hd__xnor2_2 c243 (.A(net63),
    .B(net61),
    .Y(net1008));
 sky130_fd_sc_hd__a21bo_1 c244 (.A1(net28),
    .A2(clknet_1_1__leaf_net991),
    .B1_N(net835),
    .X(net180));
 sky130_fd_sc_hd__sdfrtp_4 c245 (.CLK(clknet_4_5_0_clk),
    .D(net145),
    .RESET_B(net1002),
    .SCD(net66),
    .SCE(net150),
    .Q(net181));
 sky130_fd_sc_hd__a31o_1 c246 (.A1(net67),
    .A2(net141),
    .A3(net1021),
    .B1(clknet_1_1__leaf_net1006),
    .X(net182));
 sky130_fd_sc_hd__xnor2_1 c247 (.A(net150),
    .B(net181),
    .Y(net989));
 sky130_fd_sc_hd__a21bo_1 c248 (.A1(net61),
    .A2(net1008),
    .B1_N(net1021),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net746),
    .X(net184));
 sky130_fd_sc_hd__a31o_1 c250 (.A1(net25),
    .A2(net181),
    .A3(net898),
    .B1(clknet_1_1__leaf_net1006),
    .X(net995));
 sky130_fd_sc_hd__sdfbbn_1 c251 (.CLK_N(clknet_4_5_0_clk),
    .D(net183),
    .RESET_B(net181),
    .SCD(net981),
    .SCE(net1008),
    .SET_B(net1066),
    .Q(net186),
    .Q_N(net185));
 sky130_fd_sc_hd__a31o_1 c252 (.A1(net184),
    .A2(net181),
    .A3(net949),
    .B1(net163),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 c253 (.A(net741),
    .X(net188));
 sky130_fd_sc_hd__a21bo_1 c254 (.A1(net59),
    .A2(net185),
    .B1_N(net988),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 c255 (.A(net785),
    .X(net190));
 sky130_fd_sc_hd__a41o_1 c256 (.A1(net188),
    .A2(net63),
    .A3(net25),
    .A4(net1008),
    .B1(net981),
    .X(net1011));
 sky130_fd_sc_hd__a21bo_1 c257 (.A1(net186),
    .A2(net949),
    .B1_N(net1034),
    .X(net962));
 sky130_fd_sc_hd__a21bo_1 c258 (.A1(net190),
    .A2(net181),
    .B1_N(net962),
    .X(net968));
 sky130_fd_sc_hd__a41o_1 c259 (.A1(net180),
    .A2(net186),
    .A3(net183),
    .A4(net978),
    .B1(net1002),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net53),
    .A1(net161),
    .A2(net185),
    .A3(net162),
    .S0(net1005),
    .S1(net962),
    .X(net192));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net67),
    .A1(net1008),
    .A2(net185),
    .A3(net181),
    .S0(net1007),
    .S1(net809),
    .X(net193));
 sky130_fd_sc_hd__a41o_1 c262 (.A1(net193),
    .A2(net186),
    .A3(net61),
    .A4(net181),
    .B1(net978),
    .X(net194));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net28),
    .A1(net193),
    .A2(net60),
    .A3(clknet_1_0__leaf_net995),
    .S0(net181),
    .S1(net809),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 c264 (.A(net708),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 c265 (.A(net708),
    .X(net197));
 sky130_fd_sc_hd__buf_1 c266 (.A(net753),
    .X(net198));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net897),
    .A2(net197),
    .B1_N(net1028),
    .X(net199));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net71),
    .B(net1030),
    .Y(net200));
 sky130_fd_sc_hd__xnor2_2 c269 (.A(net196),
    .B(net1028),
    .Y(net201));
 sky130_fd_sc_hd__a21bo_1 c270 (.A1(net956),
    .A2(net201),
    .B1_N(net1033),
    .X(net202));
 sky130_fd_sc_hd__a21bo_2 c271 (.A1(net199),
    .A2(net201),
    .B1_N(net1028),
    .X(net203));
 sky130_fd_sc_hd__sdfbbp_1 c272 (.CLK(clknet_4_2_0_clk),
    .D(net1020),
    .RESET_B(net74),
    .SCD(net203),
    .SCE(net1028),
    .SET_B(net70),
    .Q(net205),
    .Q_N(net204));
 sky130_fd_sc_hd__a31o_2 c273 (.A1(net203),
    .A2(net200),
    .A3(net1020),
    .B1(net1028),
    .X(net206));
 sky130_fd_sc_hd__a31o_2 c274 (.A1(net201),
    .A2(net197),
    .A3(net899),
    .B1(net1028),
    .X(net996));
 sky130_fd_sc_hd__a31o_1 c275 (.A1(net1028),
    .A2(net897),
    .A3(net70),
    .B1(net203),
    .X(net207));
 sky130_fd_sc_hd__a21bo_1 c276 (.A1(net196),
    .A2(net996),
    .B1_N(net1030),
    .X(net208));
 sky130_fd_sc_hd__buf_1 c277 (.A(net784),
    .X(net209));
 sky130_fd_sc_hd__buf_1 c278 (.A(net755),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c279 (.A0(net209),
    .A1(net210),
    .A2(net996),
    .A3(net199),
    .S0(net1028),
    .S1(net1020),
    .X(net211));
 sky130_fd_sc_hd__sdfbbn_1 c280 (.CLK_N(clknet_4_2_0_clk),
    .D(net996),
    .RESET_B(net205),
    .SCD(net1020),
    .SCE(net211),
    .SET_B(net1030),
    .Q(net213),
    .Q_N(net212));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net213),
    .A1(net203),
    .A2(net211),
    .A3(net209),
    .S0(net200),
    .S1(net996),
    .X(net214));
 sky130_fd_sc_hd__sdfrtp_4 c282 (.CLK(clknet_4_2_0_clk),
    .D(net203),
    .RESET_B(net211),
    .SCD(net1030),
    .SCE(net807),
    .Q(net215));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(net208),
    .A1(net197),
    .A2(net996),
    .A3(net200),
    .S0(net212),
    .S1(net807),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net211),
    .A1(net213),
    .A2(net199),
    .A3(net996),
    .S0(net1020),
    .S1(net708),
    .X(net217));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net910),
    .A1(net203),
    .A2(net708),
    .A3(net733),
    .S0(net807),
    .S1(net837),
    .X(net218));
 sky130_fd_sc_hd__buf_1 c286 (.A(net755),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 c287 (.A(net755),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 c288 (.A(net753),
    .X(net221));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net941),
    .A2(net75),
    .B1_N(net1036),
    .X(net222));
 sky130_fd_sc_hd__a31o_1 c290 (.A1(net221),
    .A2(net1053),
    .A3(net1031),
    .B1(clknet_1_1__leaf_net828),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 c291 (.A(net744),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(net931),
    .A1(net86),
    .A2(net203),
    .A3(clknet_1_0__leaf_net223),
    .S0(net197),
    .S1(net1030),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net78),
    .A1(net197),
    .A2(clknet_1_0__leaf_net225),
    .A3(net224),
    .S0(clknet_1_0__leaf_net223),
    .S1(net743),
    .X(net226));
 sky130_fd_sc_hd__buf_1 c294 (.A(net761),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net219),
    .A1(clknet_1_0__leaf_net223),
    .A2(net914),
    .A3(net78),
    .S0(net1029),
    .S1(net1035),
    .X(net228));
 sky130_fd_sc_hd__buf_1 c296 (.A(net744),
    .X(net229));
 sky130_fd_sc_hd__buf_1 c297 (.A(net784),
    .X(net230));
 sky130_fd_sc_hd__a21bo_4 c298 (.A1(net70),
    .A2(net219),
    .B1_N(net914),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 c299 (.A(net1048),
    .X(net232));
 sky130_fd_sc_hd__a21bo_1 c300 (.A1(net229),
    .A2(clknet_1_0__leaf_net228),
    .B1_N(net232),
    .X(net233));
 sky130_fd_sc_hd__buf_2 c301 (.A(net755),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(net197),
    .A1(net227),
    .A2(net931),
    .A3(net927),
    .S0(net232),
    .S1(net733),
    .X(net235));
 sky130_fd_sc_hd__sdfsbp_1 c303 (.CLK(clknet_4_2_0_clk),
    .D(clknet_1_1__leaf_net233),
    .SCD(net219),
    .SCE(net234),
    .SET_B(net231),
    .Q(net237),
    .Q_N(net236));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(clknet_1_0__leaf_net225),
    .A1(net229),
    .A2(clknet_1_0__leaf_net233),
    .A3(net234),
    .S0(net205),
    .S1(net232),
    .X(net238));
 sky130_fd_sc_hd__a21bo_1 c305 (.A1(net199),
    .A2(net235),
    .B1_N(net915),
    .X(net239));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net239),
    .A2(net234),
    .A3(net237),
    .A4(net224),
    .B1(net1029),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net235),
    .A1(net231),
    .A2(net239),
    .A3(net236),
    .S0(clknet_1_1__leaf_net828),
    .S1(net838),
    .X(net241));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net213),
    .B(net921),
    .Y(net242));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net96),
    .A2(clknet_1_0__leaf_net125),
    .B1_N(net832),
    .X(net243));
 sky130_fd_sc_hd__a21bo_1 c310 (.A1(net106),
    .A2(net927),
    .B1_N(net831),
    .X(net244));
 sky130_fd_sc_hd__xnor2_2 c311 (.A(net927),
    .B(net762),
    .Y(net245));
 sky130_fd_sc_hd__xnor2_1 c312 (.A(net244),
    .B(net245),
    .Y(net246));
 sky130_fd_sc_hd__buf_1 c313 (.A(net795),
    .X(net247));
 sky130_fd_sc_hd__xnor2_1 c314 (.A(net946),
    .B(net106),
    .Y(net958));
 sky130_fd_sc_hd__clkbuf_2 c315 (.A(net783),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 c316 (.A(net747),
    .X(net249));
 sky130_fd_sc_hd__sdfsbp_1 c317 (.CLK(clknet_4_3_0_clk),
    .D(net1053),
    .SCD(clknet_1_0__leaf_net243),
    .SCE(net762),
    .SET_B(net837),
    .Q(net251),
    .Q_N(net250));
 sky130_fd_sc_hd__buf_1 c318 (.A(net777),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(clknet_1_1__leaf_net225),
    .A1(net99),
    .A2(net84),
    .A3(net942),
    .S0(net1031),
    .S1(net832),
    .X(net253));
 sky130_fd_sc_hd__xnor2_1 c320 (.A(net247),
    .B(clknet_1_1__leaf_net223),
    .Y(net254));
 sky130_fd_sc_hd__dlymetal6s2s_1 c321 (.A(net795),
    .X(net255));
 sky130_fd_sc_hd__a41o_1 c322 (.A1(net252),
    .A2(net1019),
    .A3(net247),
    .A4(net832),
    .B1(net839),
    .X(net256));
 sky130_fd_sc_hd__a31o_1 c323 (.A1(net245),
    .A2(net247),
    .A3(net231),
    .B1(net255),
    .X(net257));
 sky130_fd_sc_hd__buf_1 c324 (.A(net798),
    .X(net258));
 sky130_fd_sc_hd__sdfbbn_2 c325 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_1__leaf_net223),
    .RESET_B(clknet_1_1__leaf_net254),
    .SCD(net249),
    .SCE(net255),
    .SET_B(clknet_1_1__leaf_net243),
    .Q(net986),
    .Q_N(net259));
 sky130_fd_sc_hd__a41o_2 c326 (.A1(net249),
    .A2(net245),
    .A3(net258),
    .A4(net242),
    .B1(net837),
    .X(net260));
 sky130_fd_sc_hd__buf_2 c327 (.A(net761),
    .X(net261));
 sky130_fd_sc_hd__a31o_1 c328 (.A1(clknet_1_0__leaf_net254),
    .A2(net252),
    .A3(net261),
    .B1(net1041),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net99),
    .A1(net261),
    .A2(net212),
    .A3(clknet_1_1__leaf_net225),
    .S0(net75),
    .S1(clknet_1_0__leaf_net243),
    .X(net263));
 sky130_fd_sc_hd__sdfstp_2 c330 (.CLK(clknet_4_3_0_clk),
    .D(net942),
    .SCD(net90),
    .SCE(net155),
    .SET_B(net1064),
    .Q(net264));
 sky130_fd_sc_hd__sdfstp_1 c331 (.CLK(clknet_4_4_0_clk),
    .D(net1004),
    .SCD(net1021),
    .SCE(net155),
    .SET_B(net830),
    .Q(net265));
 sky130_fd_sc_hd__a21bo_1 c332 (.A1(net899),
    .A2(net248),
    .B1_N(net1049),
    .X(net266));
 sky130_fd_sc_hd__a21bo_2 c333 (.A1(net266),
    .A2(net151),
    .B1_N(net135),
    .X(net982));
 sky130_fd_sc_hd__sdfstp_2 c334 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net143),
    .SCD(net265),
    .SCE(net155),
    .SET_B(net1053),
    .Q(net992));
 sky130_fd_sc_hd__a21bo_1 c335 (.A1(net265),
    .A2(net248),
    .B1_N(net992),
    .X(net267));
 sky130_fd_sc_hd__a31o_1 c336 (.A1(net267),
    .A2(net982),
    .A3(net248),
    .B1(net754),
    .X(net268));
 sky130_fd_sc_hd__a41o_1 c337 (.A1(net255),
    .A2(net1019),
    .A3(clknet_1_1__leaf_net143),
    .A4(net1049),
    .B1(net942),
    .X(net269));
 sky130_fd_sc_hd__a21bo_1 c338 (.A1(net258),
    .A2(net265),
    .B1_N(net830),
    .X(net270));
 sky130_fd_sc_hd__a21bo_1 c339 (.A1(net224),
    .A2(clknet_1_0__leaf_net125),
    .B1_N(net837),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 c340 (.A(net798),
    .X(net272));
 sky130_fd_sc_hd__a31o_4 c341 (.A1(net267),
    .A2(net258),
    .A3(net224),
    .B1(net724),
    .X(net987));
 sky130_fd_sc_hd__sedfxbp_2 c342 (.CLK(clknet_4_6_0_clk),
    .D(net953),
    .DE(net987),
    .SCD(net982),
    .SCE(net724),
    .Q(net274),
    .Q_N(net273));
 sky130_fd_sc_hd__a31o_1 c343 (.A1(net120),
    .A2(net270),
    .A3(net273),
    .B1(net1031),
    .X(net275));
 sky130_fd_sc_hd__a41o_1 c344 (.A1(net270),
    .A2(net103),
    .A3(net274),
    .A4(net275),
    .B1(net248),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net276),
    .A1(net986),
    .A2(clknet_1_0__leaf_net143),
    .A3(net987),
    .S0(net151),
    .S1(net275),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net275),
    .A1(net276),
    .A2(net987),
    .A3(net982),
    .S0(net725),
    .S1(net820),
    .X(net278));
 sky130_fd_sc_hd__sdfbbp_1 c347 (.CLK(clknet_4_6_0_clk),
    .D(net232),
    .RESET_B(net273),
    .SCD(net992),
    .SCE(clknet_1_1__leaf_net243),
    .SET_B(net783),
    .Q(net280),
    .Q_N(net279));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net275),
    .A1(net135),
    .A2(net987),
    .A3(net265),
    .S0(net992),
    .S1(net783),
    .X(net281));
 sky130_fd_sc_hd__a41o_1 c349 (.A1(net281),
    .A2(net272),
    .A3(net275),
    .A4(clknet_1_1__leaf_net143),
    .B1(net725),
    .X(net282));
 sky130_fd_sc_hd__a41o_2 c350 (.A1(net135),
    .A2(net275),
    .A3(net265),
    .A4(net279),
    .B1(net826),
    .X(net283));
 sky130_fd_sc_hd__a41o_1 c351 (.A1(net283),
    .A2(net265),
    .A3(net248),
    .A4(net266),
    .B1(clknet_1_0__leaf_net984),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 c352 (.A(net798),
    .X(net285));
 sky130_fd_sc_hd__a21bo_1 c353 (.A1(net949),
    .A2(net769),
    .B1_N(clknet_1_1__leaf_net991),
    .X(net1001));
 sky130_fd_sc_hd__xnor2_1 c354 (.A(clknet_1_1__leaf_net160),
    .B(net997),
    .Y(net286));
 sky130_fd_sc_hd__a31o_1 c355 (.A1(net84),
    .A2(clknet_1_0__leaf_net271),
    .A3(net285),
    .B1(clknet_1_0__leaf_net991),
    .X(net287));
 sky130_fd_sc_hd__buf_2 c356 (.A(net760),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net141),
    .A1(net285),
    .A2(net33),
    .A3(net949),
    .S0(net288),
    .S1(net224),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c358 (.A0(net285),
    .A1(clknet_1_0__leaf_net160),
    .A2(net248),
    .A3(net288),
    .S0(net283),
    .S1(net836),
    .X(net290));
 sky130_fd_sc_hd__a21bo_1 c359 (.A1(net899),
    .A2(net167),
    .B1_N(net820),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 c360 (.A(net785),
    .X(net292));
 sky130_fd_sc_hd__a21bo_1 c361 (.A1(net175),
    .A2(net1004),
    .B1_N(net288),
    .X(net975));
 sky130_fd_sc_hd__a21bo_1 c362 (.A1(net174),
    .A2(net288),
    .B1_N(net833),
    .X(net293));
 sky130_fd_sc_hd__a31o_1 c363 (.A1(net292),
    .A2(net175),
    .A3(net1034),
    .B1(net1013),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 c364 (.A(net784),
    .X(net295));
 sky130_fd_sc_hd__buf_1 c365 (.A(net798),
    .X(net296));
 sky130_fd_sc_hd__a21bo_2 c366 (.A1(net248),
    .A2(net975),
    .B1_N(net997),
    .X(net983));
 sky130_fd_sc_hd__a21bo_1 c367 (.A1(net167),
    .A2(net215),
    .B1_N(net820),
    .X(net297));
 sky130_fd_sc_hd__a21bo_1 c368 (.A1(net295),
    .A2(net710),
    .B1_N(net811),
    .X(net298));
 sky130_fd_sc_hd__a21bo_1 c369 (.A1(net298),
    .A2(net141),
    .B1_N(net754),
    .X(net299));
 sky130_fd_sc_hd__a21bo_1 c370 (.A1(net296),
    .A2(net297),
    .B1_N(net997),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_1 c371 (.A(net784),
    .X(net300));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net299),
    .A1(net292),
    .A2(net300),
    .A3(net288),
    .S0(net1045),
    .S1(clknet_1_0__leaf_net1001),
    .X(net973));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net300),
    .A1(net283),
    .A2(net167),
    .A3(net179),
    .S0(net296),
    .S1(net987),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net283),
    .A1(clknet_1_0__leaf_net973),
    .A2(net1004),
    .A3(net141),
    .S0(clknet_1_0__leaf_net995),
    .S1(net811),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net291),
    .A1(net295),
    .A2(net983),
    .A3(net1004),
    .S0(net998),
    .S1(net840),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net162),
    .A1(net1019),
    .A2(net809),
    .A3(net997),
    .S0(net1091),
    .S1(net1075),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net161),
    .A1(net195),
    .A2(net1005),
    .S0(net964),
    .S1(net841),
    .X(net305));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net92),
    .B(net86),
    .Y(net306));
 sky130_fd_sc_hd__xnor2_2 c397 (.A(net907),
    .B(net306),
    .Y(net307));
 sky130_fd_sc_hd__clkbuf_2 c398 (.A(net717),
    .X(net308));
 sky130_fd_sc_hd__buf_1 c399 (.A(net717),
    .X(net309));
 sky130_fd_sc_hd__a31o_4 c400 (.A1(net306),
    .A2(net952),
    .A3(net308),
    .B1(net1028),
    .X(net310));
 sky130_fd_sc_hd__buf_2 c401 (.A(net663),
    .X(net311));
 sky130_fd_sc_hd__xnor2_1 c402 (.A(net1022),
    .B(net306),
    .Y(net312));
 sky130_fd_sc_hd__a21bo_1 c403 (.A1(net955),
    .A2(net85),
    .B1_N(net311),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_2 c404 (.A(net717),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 c405 (.A(net670),
    .X(net314));
 sky130_fd_sc_hd__a41o_2 c406 (.A1(net314),
    .A2(net313),
    .A3(net308),
    .A4(net196),
    .B1(net1033),
    .X(net315));
 sky130_fd_sc_hd__xnor2_2 c407 (.A(net313),
    .B(net1018),
    .Y(net316));
 sky130_fd_sc_hd__buf_6 c408 (.A(net775),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 c409 (.A(net670),
    .X(net318));
 sky130_fd_sc_hd__xnor2_4 c410 (.A(net306),
    .B(net318),
    .Y(net319));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(net308),
    .A2(net316),
    .B1_N(net313),
    .X(net320));
 sky130_fd_sc_hd__xnor2_1 c412 (.A(net315),
    .B(net319),
    .Y(net321));
 sky130_fd_sc_hd__buf_1 c413 (.A(net790),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 c414 (.A(net815),
    .X(net323));
 sky130_fd_sc_hd__xnor2_2 c415 (.A(net908),
    .B(net910),
    .Y(net324));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net320),
    .A1(net324),
    .A2(net323),
    .A3(net313),
    .S0(net1022),
    .S1(net1028),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net210),
    .A1(net310),
    .A2(net323),
    .A3(net89),
    .S0(net320),
    .S1(net842),
    .X(net326));
 sky130_fd_sc_hd__buf_2 c418 (.A(net719),
    .X(net327));
 sky130_fd_sc_hd__buf_1 c419 (.A(net718),
    .X(net328));
 sky130_fd_sc_hd__a21bo_2 c420 (.A1(net323),
    .A2(net956),
    .B1_N(net230),
    .X(net1010));
 sky130_fd_sc_hd__a21bo_1 c421 (.A1(net227),
    .A2(net234),
    .B1_N(net328),
    .X(net329));
 sky130_fd_sc_hd__a21bo_1 c422 (.A1(net203),
    .A2(net1036),
    .B1_N(net196),
    .X(net330));
 sky130_fd_sc_hd__a21bo_1 c423 (.A1(net329),
    .A2(net110),
    .B1_N(net227),
    .X(net331));
 sky130_fd_sc_hd__buf_1 c424 (.A(net719),
    .X(net332));
 sky130_fd_sc_hd__xnor2_1 c425 (.A(net110),
    .B(net842),
    .Y(net333));
 sky130_fd_sc_hd__xnor2_1 c426 (.A(net333),
    .B(net313),
    .Y(net334));
 sky130_fd_sc_hd__a21bo_1 c427 (.A1(net328),
    .A2(net332),
    .B1_N(net322),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(net316),
    .A1(net330),
    .A2(net333),
    .A3(net206),
    .S0(net327),
    .S1(net1038),
    .X(net336));
 sky130_fd_sc_hd__a21bo_1 c429 (.A1(net334),
    .A2(net327),
    .B1_N(net844),
    .X(net337));
 sky130_fd_sc_hd__a21bo_1 c430 (.A1(net220),
    .A2(net316),
    .B1_N(net844),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net313),
    .A1(net1020),
    .A2(net332),
    .A3(net338),
    .S0(net327),
    .S1(net331),
    .X(net339));
 sky130_fd_sc_hd__a21bo_2 c432 (.A1(net955),
    .A2(net96),
    .B1_N(net844),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net206),
    .A1(net1018),
    .A2(net329),
    .A3(net316),
    .S0(net332),
    .S1(net327),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 c434 (.A(net718),
    .X(net342));
 sky130_fd_sc_hd__a21bo_1 c435 (.A1(net220),
    .A2(net323),
    .B1_N(clknet_1_0__leaf_net845),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net332),
    .A1(net338),
    .A2(net342),
    .A3(net89),
    .S0(net335),
    .S1(clknet_1_0__leaf_net845),
    .X(net344));
 sky130_fd_sc_hd__buf_1 c437 (.A(net717),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net343),
    .A1(net320),
    .A2(net918),
    .A3(net1020),
    .S0(net316),
    .S1(clknet_1_0__leaf_net847),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net335),
    .A1(net329),
    .A2(net328),
    .A3(net322),
    .S0(net842),
    .S1(net848),
    .X(net347));
 sky130_fd_sc_hd__sedfxbp_1 c440 (.CLK(clknet_4_3_0_clk),
    .D(net262),
    .DE(net331),
    .SCD(net812),
    .SCE(net1042),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__buf_1 c441 (.A(clknet_1_0__leaf_net792),
    .X(net350));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net327),
    .A2(net308),
    .B1_N(net348),
    .X(net351));
 sky130_fd_sc_hd__xnor2_1 c443 (.A(net261),
    .B(net310),
    .Y(net352));
 sky130_fd_sc_hd__xnor2_1 c444 (.A(clknet_1_0__leaf_net350),
    .B(net92),
    .Y(net353));
 sky130_fd_sc_hd__a31o_1 c445 (.A1(net318),
    .A2(clknet_1_0__leaf_net353),
    .A3(net351),
    .B1(net260),
    .X(net354));
 sky130_fd_sc_hd__buf_1 c446 (.A(clknet_1_0__leaf_net792),
    .X(net355));
 sky130_fd_sc_hd__buf_1 c447 (.A(net963),
    .X(net356));
 sky130_fd_sc_hd__xnor2_1 c448 (.A(net331),
    .B(clknet_1_1__leaf_net353),
    .Y(net357));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net356),
    .A1(net901),
    .A2(clknet_1_1__leaf_net350),
    .A3(net318),
    .S0(net1042),
    .S1(clknet_1_0__leaf_net847),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 c450 (.A(net789),
    .X(net359));
 sky130_fd_sc_hd__a41o_1 c451 (.A1(net230),
    .A2(clknet_1_1__leaf_net353),
    .A3(clknet_1_0__leaf_net357),
    .A4(net345),
    .B1(net356),
    .X(net360));
 sky130_fd_sc_hd__xnor2_4 c452 (.A(net310),
    .B(net260),
    .Y(net361));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(clknet_1_1__leaf_net355),
    .A1(net327),
    .A2(net947),
    .A3(net261),
    .S0(net1015),
    .S1(clknet_1_1__leaf_net353),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 c454 (.A(net744),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(net352),
    .A1(net308),
    .A2(net337),
    .A3(net327),
    .S0(net1015),
    .S1(net318),
    .X(net364));
 sky130_fd_sc_hd__sedfxtp_4 c456 (.CLK(clknet_4_12_0_clk),
    .D(net927),
    .DE(net351),
    .SCD(net1015),
    .SCE(net812),
    .Q(net969));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net256),
    .A1(net123),
    .A2(clknet_1_0__leaf_net353),
    .A3(net349),
    .S0(net261),
    .S1(net852),
    .X(net365));
 sky130_fd_sc_hd__sdfbbn_1 c458 (.CLK_N(clknet_4_9_0_clk),
    .D(net260),
    .RESET_B(net1016),
    .SCD(net1040),
    .SCE(net853),
    .SET_B(net1069),
    .Q(net367),
    .Q_N(net366));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net367),
    .A1(net1092),
    .A2(net310),
    .A3(net318),
    .S0(net1015),
    .S1(net1067),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net261),
    .A1(net366),
    .A2(net969),
    .A3(net1016),
    .S0(net716),
    .S1(net854),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(clknet_1_1__leaf_net358),
    .A1(net366),
    .A2(net330),
    .A3(net318),
    .S0(net716),
    .S1(net853),
    .X(net370));
 sky130_fd_sc_hd__a31o_1 c462 (.A1(net215),
    .A2(net1018),
    .A3(net1017),
    .B1(net716),
    .X(net371));
 sky130_fd_sc_hd__a31o_1 c463 (.A1(net151),
    .A2(net986),
    .A3(net1031),
    .B1(net1015),
    .X(net372));
 sky130_fd_sc_hd__a21bo_1 c464 (.A1(net1022),
    .A2(net280),
    .B1_N(net151),
    .X(net373));
 sky130_fd_sc_hd__a21bo_1 c465 (.A1(net135),
    .A2(net232),
    .B1_N(clknet_1_0__leaf_net793),
    .X(net374));
 sky130_fd_sc_hd__a21bo_1 c466 (.A1(net751),
    .A2(clknet_1_0__leaf_net793),
    .B1_N(net800),
    .X(net971));
 sky130_fd_sc_hd__a31o_1 c467 (.A1(net921),
    .A2(clknet_1_0__leaf_net119),
    .A3(net1017),
    .B1(net785),
    .X(net375));
 sky130_fd_sc_hd__a21bo_1 c468 (.A1(net1045),
    .A2(net1018),
    .B1_N(net953),
    .X(net376));
 sky130_fd_sc_hd__buf_1 c469 (.A(net797),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 c470 (.A(net797),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_1 c471 (.A(net804),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net378),
    .A1(net351),
    .A2(clknet_1_0__leaf_net971),
    .A3(net264),
    .S0(net785),
    .S1(net854),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net1031),
    .A1(clknet_1_0__leaf_net379),
    .A2(net377),
    .A3(net1018),
    .S0(net987),
    .S1(net751),
    .X(net380));
 sky130_fd_sc_hd__a21bo_1 c474 (.A1(net351),
    .A2(clknet_1_0__leaf_net971),
    .B1_N(net716),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 c475 (.A(net804),
    .X(net967));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(clknet_1_0__leaf_net380),
    .A1(net953),
    .A2(net1027),
    .A3(net1026),
    .S0(net1015),
    .S1(net1031),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net232),
    .A1(net378),
    .A2(clknet_1_0__leaf_net380),
    .A3(clknet_1_0__leaf_net381),
    .S0(net1018),
    .S1(net1031),
    .X(net383));
 sky130_fd_sc_hd__a31o_1 c478 (.A1(clknet_1_0__leaf_net380),
    .A2(net1018),
    .A3(net1026),
    .B1(net747),
    .X(net384));
 sky130_fd_sc_hd__a31o_1 c479 (.A1(net345),
    .A2(net1027),
    .A3(clknet_1_0__leaf_net379),
    .B1(net1026),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net385),
    .A1(net377),
    .A2(net151),
    .A3(net953),
    .S0(net272),
    .S1(clknet_1_0__leaf_net381),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net377),
    .A1(clknet_1_1__leaf_net380),
    .A2(clknet_1_0__leaf_net379),
    .A3(net272),
    .S0(net803),
    .S1(net814),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net380),
    .A1(clknet_1_0__leaf_net379),
    .A2(net232),
    .A3(net376),
    .S0(net814),
    .S1(net854),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net1018),
    .A1(net232),
    .A2(clknet_1_0__leaf_net971),
    .A3(net791),
    .S0(net803),
    .S1(net855),
    .X(net389));
 sky130_fd_sc_hd__a41o_1 c484 (.A1(net1021),
    .A2(net1034),
    .A3(clknet_1_0__leaf_net286),
    .A4(net288),
    .B1(net836),
    .X(net976));
 sky130_fd_sc_hd__sedfxtp_4 c485 (.CLK(clknet_4_6_0_clk),
    .D(net89),
    .DE(net969),
    .SCD(net1045),
    .SCE(net834),
    .Q(net390));
 sky130_fd_sc_hd__a41o_1 c486 (.A1(net960),
    .A2(net983),
    .A3(clknet_1_1__leaf_net125),
    .A4(net800),
    .B1(net836),
    .X(net391));
 sky130_fd_sc_hd__sedfxtp_2 c487 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net125),
    .DE(net974),
    .SCD(net1018),
    .SCE(net960),
    .Q(net392));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net392),
    .A1(net1013),
    .A2(net1019),
    .A3(net373),
    .S0(clknet_1_1__leaf_net792),
    .S1(net794),
    .X(net393));
 sky130_fd_sc_hd__sdfbbn_1 c489 (.CLK_N(clknet_4_6_0_clk),
    .D(net373),
    .RESET_B(net215),
    .SCD(net1027),
    .SCE(net259),
    .SET_B(net915),
    .Q(net972),
    .Q_N(net394));
 sky130_fd_sc_hd__sdfrbp_1 c490 (.CLK(clknet_4_7_0_clk),
    .D(net179),
    .RESET_B(clknet_1_0__leaf_net164),
    .SCD(net972),
    .SCE(net983),
    .Q(net396),
    .Q_N(net395));
 sky130_fd_sc_hd__a41o_1 c491 (.A1(net396),
    .A2(clknet_1_1__leaf_net125),
    .A3(net33),
    .A4(net392),
    .B1(net814),
    .X(net397));
 sky130_fd_sc_hd__a41o_1 c492 (.A1(net901),
    .A2(net975),
    .A3(net974),
    .A4(net394),
    .B1(clknet_1_1__leaf_net846),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_1__leaf_net966),
    .A1(net394),
    .A2(net288),
    .A3(clknet_1_1__leaf_net750),
    .S0(net813),
    .S1(clknet_1_0__leaf_net991),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net398),
    .A1(net1026),
    .A2(net293),
    .A3(net394),
    .S0(clknet_1_0__leaf_net164),
    .S1(clknet_1_0__leaf_net991),
    .X(net400));
 sky130_fd_sc_hd__a41o_1 c495 (.A1(net902),
    .A2(net395),
    .A3(net390),
    .A4(clknet_1_1__leaf_net792),
    .B1(net856),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net390),
    .A1(net396),
    .A2(net921),
    .A3(net1027),
    .S0(clknet_1_0__leaf_net971),
    .S1(clknet_1_1__leaf_net846),
    .X(net402));
 sky130_fd_sc_hd__a41o_1 c497 (.A1(net972),
    .A2(net33),
    .A3(net1027),
    .A4(net759),
    .B1(net836),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net215),
    .A1(net1036),
    .A2(net972),
    .A3(clknet_1_1__leaf_net750),
    .S0(clknet_1_0__leaf_net984),
    .S1(net856),
    .X(net404));
 sky130_fd_sc_hd__a41o_1 c499 (.A1(net396),
    .A2(net178),
    .A3(net979),
    .A4(clknet_1_1__leaf_net846),
    .B1(net856),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(clknet_1_0__leaf_net405),
    .A1(net33),
    .A2(clknet_1_0__leaf_net404),
    .A3(net1017),
    .S0(clknet_1_0__leaf_net991),
    .S1(net1073),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net288),
    .A1(clknet_1_0__leaf_net404),
    .A2(net1034),
    .A3(net993),
    .S0(net836),
    .S1(net857),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(clknet_1_0__leaf_net407),
    .A1(net914),
    .A2(clknet_1_0__leaf_net404),
    .A3(net178),
    .S0(net395),
    .S1(net856),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net392),
    .A1(clknet_1_0__leaf_net404),
    .A2(clknet_1_1__leaf_net405),
    .A3(net993),
    .S0(net839),
    .S1(net857),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net401),
    .A1(net288),
    .A2(clknet_1_1__leaf_net407),
    .A3(net390),
    .S0(clknet_1_0__leaf_net409),
    .S1(net1050),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net408),
    .A1(clknet_1_0__leaf_net407),
    .A2(net1013),
    .A3(net392),
    .S0(net1026),
    .S1(net759),
    .X(net411));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net76),
    .B(net1038),
    .Y(net412));
 sky130_fd_sc_hd__buf_2 c529 (.A(net712),
    .X(net413));
 sky130_fd_sc_hd__xnor2_2 c530 (.A(net910),
    .B(net314),
    .Y(net414));
 sky130_fd_sc_hd__xnor2_4 c531 (.A(net319),
    .B(net412),
    .Y(net415));
 sky130_fd_sc_hd__buf_1 c532 (.A(net711),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 c533 (.A(net682),
    .X(net417));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net311),
    .B(net76),
    .Y(net418));
 sky130_fd_sc_hd__mux4_1 c535 (.A0(net904),
    .A1(net311),
    .A2(net315),
    .A3(net418),
    .S0(net415),
    .S1(net412),
    .X(net419));
 sky130_fd_sc_hd__xnor2_2 c536 (.A(net314),
    .B(net1040),
    .Y(net420));
 sky130_fd_sc_hd__clkbuf_2 c537 (.A(net681),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net417),
    .A1(net420),
    .A2(net317),
    .A3(net412),
    .S0(net415),
    .S1(net413),
    .X(net422));
 sky130_fd_sc_hd__a21bo_1 c539 (.A1(net309),
    .A2(net416),
    .B1_N(net862),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 c540 (.A(net790),
    .X(net424));
 sky130_fd_sc_hd__a21bo_4 c541 (.A1(net317),
    .A2(net311),
    .B1_N(net1088),
    .X(net425));
 sky130_fd_sc_hd__a41o_1 c542 (.A1(net414),
    .A2(net421),
    .A3(net416),
    .A4(net218),
    .B1(net76),
    .X(net426));
 sky130_fd_sc_hd__buf_1 c543 (.A(net700),
    .X(net427));
 sky130_fd_sc_hd__a21bo_1 c544 (.A1(net427),
    .A2(net1024),
    .B1_N(net860),
    .X(net428));
 sky130_fd_sc_hd__a41o_2 c545 (.A1(net412),
    .A2(net418),
    .A3(net427),
    .A4(net1024),
    .B1(net859),
    .X(net429));
 sky130_fd_sc_hd__xnor2_2 c546 (.A(net423),
    .B(net428),
    .Y(net430));
 sky130_fd_sc_hd__mux4_2 c547 (.A0(net428),
    .A1(net430),
    .A2(net429),
    .A3(net421),
    .S0(net423),
    .S1(net311),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 c548 (.A(net699),
    .X(net432));
 sky130_fd_sc_hd__mux4_2 c549 (.A0(net432),
    .A1(net427),
    .A2(net412),
    .A3(net309),
    .S0(net712),
    .S1(net860),
    .X(net433));
 sky130_fd_sc_hd__xnor2_4 c550 (.A(net429),
    .B(net1047),
    .Y(net434));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net901),
    .A2(net1010),
    .B1_N(net896),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 c552 (.A(net732),
    .X(net436));
 sky130_fd_sc_hd__sdfrbp_1 c553 (.CLK(clknet_4_8_0_clk),
    .D(net324),
    .RESET_B(net342),
    .SCD(net1010),
    .SCE(net434),
    .Q(net438),
    .Q_N(net437));
 sky130_fd_sc_hd__a21bo_1 c554 (.A1(net436),
    .A2(net429),
    .B1_N(net1020),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 c555 (.A(net731),
    .X(net440));
 sky130_fd_sc_hd__buf_1 c556 (.A(net1074),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(net435),
    .A1(net1010),
    .A2(net434),
    .A3(net202),
    .S0(net1033),
    .S1(clknet_1_1__leaf_net847),
    .X(net442));
 sky130_fd_sc_hd__buf_1 c558 (.A(net742),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net732),
    .X(net444));
 sky130_fd_sc_hd__xnor2_2 c560 (.A(net421),
    .B(net863),
    .Y(net445));
 sky130_fd_sc_hd__a21bo_1 c561 (.A1(net435),
    .A2(net443),
    .B1_N(net440),
    .X(net446));
 sky130_fd_sc_hd__sdfbbp_1 c562 (.CLK(clknet_4_9_0_clk),
    .D(net443),
    .RESET_B(net340),
    .SCD(net96),
    .SCE(net439),
    .SET_B(net441),
    .Q(net448),
    .Q_N(net447));
 sky130_fd_sc_hd__buf_2 c563 (.A(net742),
    .X(net999));
 sky130_fd_sc_hd__dlymetal6s2s_1 c564 (.A(net744),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net438),
    .A1(net338),
    .A2(net449),
    .A3(net436),
    .S0(net342),
    .S1(net234),
    .X(net450));
 sky130_fd_sc_hd__a21bo_1 c566 (.A1(clknet_1_1__leaf_net845),
    .A2(net863),
    .B1_N(net864),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_0__leaf_net451),
    .A1(net430),
    .A2(net420),
    .A3(net110),
    .S0(net236),
    .S1(net1047),
    .X(net452));
 sky130_fd_sc_hd__a21bo_1 c568 (.A1(net956),
    .A2(net440),
    .B1_N(net864),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net896),
    .A1(net999),
    .A2(clknet_1_0__leaf_net452),
    .A3(net443),
    .S0(net447),
    .S1(net864),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net449),
    .A1(net453),
    .A2(net1022),
    .A3(clknet_1_1__leaf_net451),
    .S0(net443),
    .S1(net437),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net453),
    .A1(net445),
    .A2(net444),
    .A3(net438),
    .S0(clknet_1_0__leaf_net455),
    .S1(net864),
    .X(net456));
 sky130_fd_sc_hd__a21bo_1 c572 (.A1(net96),
    .A2(net413),
    .B1_N(net1033),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 c573 (.A(net791),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(net453),
    .A1(net359),
    .A2(net441),
    .A3(net434),
    .S0(net812),
    .S1(net1040),
    .X(net459));
 sky130_fd_sc_hd__xnor2_1 c575 (.A(net367),
    .B(net449),
    .Y(net460));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net791),
    .X(net461));
 sky130_fd_sc_hd__buf_1 c577 (.A(clknet_1_0__leaf_net749),
    .X(net462));
 sky130_fd_sc_hd__buf_1 c578 (.A(net789),
    .X(net463));
 sky130_fd_sc_hd__xnor2_1 c579 (.A(net941),
    .B(net433),
    .Y(net464));
 sky130_fd_sc_hd__buf_1 c580 (.A(clknet_1_1__leaf_net662),
    .X(net465));
 sky130_fd_sc_hd__a21bo_1 c581 (.A1(net465),
    .A2(net969),
    .B1_N(net250),
    .X(net466));
 sky130_fd_sc_hd__buf_1 c582 (.A(net742),
    .X(net467));
 sky130_fd_sc_hd__a21bo_1 c583 (.A1(net441),
    .A2(net463),
    .B1_N(net1040),
    .X(net468));
 sky130_fd_sc_hd__a31o_1 c584 (.A1(net363),
    .A2(net1024),
    .A3(net440),
    .B1(net1032),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net466),
    .A1(net337),
    .A2(net433),
    .A3(net440),
    .S0(net1015),
    .S1(net1032),
    .X(net470));
 sky130_fd_sc_hd__xnor2_1 c586 (.A(net251),
    .B(clknet_1_1__leaf_net119),
    .Y(net471));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(net468),
    .A1(clknet_1_0__leaf_net455),
    .A2(net440),
    .A3(net1016),
    .S0(clknet_1_0__leaf_net847),
    .S1(net851),
    .X(net472));
 sky130_fd_sc_hd__a21bo_1 c588 (.A1(net251),
    .A2(clknet_1_1__leaf_net749),
    .B1_N(clknet_1_0__leaf_net867),
    .X(net959));
 sky130_fd_sc_hd__buf_1 c589 (.A(clknet_1_0__leaf_net662),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net471),
    .A1(net473),
    .A2(net441),
    .A3(net467),
    .S0(net434),
    .S1(net433),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net462),
    .A1(net469),
    .A2(net340),
    .A3(net1024),
    .S0(net1040),
    .S1(clknet_1_0__leaf_net847),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net460),
    .A1(net463),
    .A2(net851),
    .A3(clknet_1_0__leaf_net867),
    .S0(clknet_1_0__leaf_net961),
    .S1(net869),
    .X(net476));
 sky130_fd_sc_hd__a21bo_1 c593 (.A1(clknet_1_1__leaf_net867),
    .A2(clknet_1_0__leaf_net961),
    .B1_N(net869),
    .X(net477));
 sky130_fd_sc_hd__sdfbbn_1 c594 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net455),
    .RESET_B(net1049),
    .SCD(net274),
    .SCE(net1019),
    .SET_B(clknet_1_1__leaf_net381),
    .Q(net479),
    .Q_N(net478));
 sky130_fd_sc_hd__a41o_1 c595 (.A1(net272),
    .A2(clknet_1_0__leaf_net476),
    .A3(clknet_1_1__leaf_net381),
    .A4(net89),
    .B1(net1045),
    .X(net480));
 sky130_fd_sc_hd__sdfbbn_1 c596 (.CLK_N(clknet_4_12_0_clk),
    .D(net446),
    .RESET_B(net448),
    .SCD(clknet_1_0__leaf_net452),
    .SCE(net1015),
    .SET_B(net1032),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__sdfbbp_1 c597 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net389),
    .RESET_B(net479),
    .SCD(clknet_1_1__leaf_net966),
    .SCE(net1024),
    .SET_B(net1085),
    .Q(net484),
    .Q_N(net483));
 sky130_fd_sc_hd__sdfrtn_1 c598 (.CLK_N(clknet_4_11_0_clk),
    .D(net359),
    .RESET_B(net1016),
    .SCD(net440),
    .SCE(net447),
    .Q(net485));
 sky130_fd_sc_hd__sdfbbn_1 c599 (.CLK_N(clknet_4_12_0_clk),
    .D(net446),
    .RESET_B(net969),
    .SCD(net413),
    .SCE(net376),
    .SET_B(net1042),
    .Q(net487),
    .Q_N(net486));
 sky130_fd_sc_hd__mux4_2 c600 (.A0(net482),
    .A1(net483),
    .A2(net274),
    .A3(net486),
    .S0(net1032),
    .S1(net901),
    .X(net488));
 sky130_fd_sc_hd__sdfbbn_2 c601 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net455),
    .RESET_B(net1024),
    .SCD(net791),
    .SCE(net833),
    .SET_B(net1065),
    .Q(net490),
    .Q_N(net489));
 sky130_fd_sc_hd__a41o_1 c602 (.A1(net440),
    .A2(clknet_1_0__leaf_net476),
    .A3(net1024),
    .A4(net481),
    .B1(clknet_1_0__leaf_net846),
    .X(net491));
 sky130_fd_sc_hd__a41o_1 c603 (.A1(net376),
    .A2(net487),
    .A3(net280),
    .A4(net819),
    .B1(net833),
    .X(net492));
 sky130_fd_sc_hd__a41o_1 c604 (.A1(net434),
    .A2(net482),
    .A3(net488),
    .A4(clknet_1_1__leaf_net389),
    .B1(net1026),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_1__leaf_net381),
    .A1(net999),
    .A2(net481),
    .A3(net1037),
    .S0(net446),
    .S1(net273),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net918),
    .A1(clknet_1_0__leaf_net491),
    .A2(net1016),
    .A3(net801),
    .S0(net1042),
    .S1(net990),
    .X(net495));
 sky130_fd_sc_hd__a41o_1 c607 (.A1(clknet_1_1__leaf_net379),
    .A2(net1027),
    .A3(net1042),
    .A4(net849),
    .B1(net990),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net484),
    .A1(clknet_1_1__leaf_net452),
    .A2(net1022),
    .A3(clknet_1_1__leaf_net379),
    .S0(net481),
    .S1(net870),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(net496),
    .A1(clknet_1_0__leaf_net491),
    .A2(clknet_1_1__leaf_net379),
    .A3(net868),
    .S0(net870),
    .S1(net871),
    .X(net498));
 sky130_fd_sc_hd__a41o_1 c610 (.A1(net274),
    .A2(net482),
    .A3(net486),
    .A4(net834),
    .B1(net871),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net488),
    .A1(net489),
    .A2(net801),
    .A3(clknet_1_1__leaf_net867),
    .S0(net990),
    .S1(net872),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(clknet_1_0__leaf_net500),
    .A1(net484),
    .A2(net1037),
    .A3(net479),
    .S0(net1026),
    .S1(net870),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net499),
    .A1(clknet_1_1__leaf_net501),
    .A2(net1024),
    .A3(clknet_1_1__leaf_net500),
    .S0(net376),
    .S1(net819),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(clknet_1_0__leaf_net501),
    .A1(clknet_1_0__leaf_net500),
    .A2(net478),
    .A3(net279),
    .S0(net808),
    .S1(net872),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net340),
    .A1(net492),
    .A2(net1044),
    .A3(net1017),
    .S0(clknet_1_0__leaf_net501),
    .S1(net488),
    .X(net504));
 sky130_fd_sc_hd__sdfbbp_1 c616 (.CLK(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net404),
    .RESET_B(net1024),
    .SCD(net1034),
    .SCE(clknet_1_1__leaf_net966),
    .SET_B(net1026),
    .Q(net506),
    .Q_N(net505));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net464),
    .A1(net390),
    .A2(net488),
    .A3(net921),
    .S0(net1027),
    .S1(net905),
    .X(net507));
 sky130_fd_sc_hd__a41o_1 c618 (.A1(net402),
    .A2(net424),
    .A3(net490),
    .A4(clknet_1_1__leaf_net164),
    .B1(net279),
    .X(net508));
 sky130_fd_sc_hd__a41o_1 c619 (.A1(net280),
    .A2(net506),
    .A3(net1027),
    .A4(net488),
    .B1(net858),
    .X(net509));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net937),
    .A1(net942),
    .A2(net948),
    .A3(net944),
    .S0(net940),
    .S1(net911),
    .X(net0));
 sky130_fd_sc_hd__sdfbbn_1 c620 (.CLK_N(clknet_4_13_0_clk),
    .D(net509),
    .RESET_B(clknet_1_1__leaf_net476),
    .SCD(net922),
    .SCE(clknet_1_1__leaf_net164),
    .SET_B(net505),
    .Q(net511),
    .Q_N(net510));
 sky130_fd_sc_hd__a41o_1 c621 (.A1(net488),
    .A2(net1019),
    .A3(net33),
    .A4(net707),
    .B1(net1050),
    .X(net512));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net511),
    .A1(clknet_1_1__leaf_net164),
    .A2(net1027),
    .A3(net1009),
    .S0(clknet_1_1__leaf_net749),
    .S1(net802),
    .X(net513));
 sky130_fd_sc_hd__a41o_1 c623 (.A1(net511),
    .A2(net909),
    .A3(net424),
    .A4(clknet_1_1__leaf_net164),
    .B1(net1017),
    .X(net514));
 sky130_fd_sc_hd__a41o_1 c624 (.A1(net921),
    .A2(net1027),
    .A3(net1026),
    .A4(net772),
    .B1(net855),
    .X(net515));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(clknet_1_1__leaf_net164),
    .A1(net390),
    .A2(net999),
    .A3(net921),
    .S0(net510),
    .S1(net858),
    .X(net516));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(clknet_1_1__leaf_net286),
    .A1(net453),
    .A2(net506),
    .A3(net489),
    .S0(clknet_1_1__leaf_net164),
    .S1(net980),
    .X(net517));
 sky130_fd_sc_hd__a41o_1 c627 (.A1(net33),
    .A2(net488),
    .A3(net970),
    .A4(net1082),
    .B1(net980),
    .X(net518));
 sky130_fd_sc_hd__a41o_1 c628 (.A1(net921),
    .A2(net485),
    .A3(clknet_1_1__leaf_net404),
    .A4(net707),
    .B1(net874),
    .X(net519));
 sky130_fd_sc_hd__a41o_1 c629 (.A1(net1089),
    .A2(net515),
    .A3(net33),
    .A4(net980),
    .B1(net874),
    .X(net520));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net924),
    .A1(net945),
    .A2(net944),
    .A3(net950),
    .S0(net946),
    .S1(net911),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net293),
    .A1(clknet_1_1__leaf_net404),
    .A2(net1045),
    .A3(net1017),
    .S0(net977),
    .S1(net980),
    .X(net521));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net461),
    .A1(net983),
    .A2(net1017),
    .A3(net813),
    .S0(net980),
    .S1(net1086),
    .X(net522));
 sky130_fd_sc_hd__a41o_1 c632 (.A1(clknet_1_1__leaf_net971),
    .A2(net772),
    .A3(net980),
    .A4(net874),
    .B1(net875),
    .X(net523));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(clknet_1_1__leaf_net357),
    .A1(net509),
    .A2(clknet_1_1__leaf_net404),
    .A3(net858),
    .S0(net980),
    .S1(net875),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net523),
    .A1(clknet_1_1__leaf_net971),
    .A2(net390),
    .A3(net758),
    .S0(net980),
    .S1(net875),
    .X(net525));
 sky130_fd_sc_hd__a41o_1 c635 (.A1(net525),
    .A2(net857),
    .A3(net980),
    .A4(net874),
    .B1(net875),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net519),
    .A1(clknet_1_0__leaf_net409),
    .A2(net1013),
    .A3(clknet_1_1__leaf_net793),
    .S0(net858),
    .S1(net875),
    .X(net527));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_4_13_0_clk),
    .D(clknet_1_1__leaf_net452),
    .RESET_B(net1010),
    .SCD(clknet_1_1__leaf_net793),
    .SCE(net875),
    .SET_B(net876),
    .Q(net529),
    .Q_N(net528));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net938),
    .A1(net1),
    .A2(net936),
    .A3(net939),
    .S0(net3),
    .S1(net947),
    .X(net2));
 sky130_fd_sc_hd__a21bo_1 c65 (.A1(net911),
    .A2(net957),
    .B1_N(net924),
    .X(net3));
 sky130_fd_sc_hd__xnor2_2 c66 (.A(net0),
    .B(net935),
    .Y(net4));
 sky130_fd_sc_hd__xnor2_2 c660 (.A(net1038),
    .B(net315),
    .Y(net530));
 sky130_fd_sc_hd__a31o_1 c661 (.A1(net315),
    .A2(net430),
    .A3(net431),
    .B1(net1088),
    .X(net531));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net530),
    .B(net414),
    .Y(net532));
 sky130_fd_sc_hd__clkbuf_1 c663 (.A(net782),
    .X(net533));
 sky130_fd_sc_hd__buf_1 c664 (.A(net782),
    .X(net534));
 sky130_fd_sc_hd__xnor2_1 c665 (.A(net904),
    .B(net1070),
    .Y(net535));
 sky130_fd_sc_hd__sdfrtp_2 c666 (.CLK(clknet_4_10_0_clk),
    .D(net532),
    .RESET_B(net534),
    .SCD(net715),
    .SCE(net1040),
    .Q(net536));
 sky130_fd_sc_hd__clkbuf_1 c667 (.A(net816),
    .X(net537));
 sky130_fd_sc_hd__xnor2_4 c668 (.A(net425),
    .B(net534),
    .Y(net538));
 sky130_fd_sc_hd__xnor2_2 c669 (.A(net538),
    .B(net862),
    .Y(net539));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net908),
    .B(net955),
    .Y(net5));
 sky130_fd_sc_hd__xnor2_1 c670 (.A(net536),
    .B(net862),
    .Y(net540));
 sky130_fd_sc_hd__buf_2 c671 (.A(net663),
    .X(net541));
 sky130_fd_sc_hd__xnor2_1 c672 (.A(net541),
    .B(net1040),
    .Y(net542));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(net210),
    .A1(net431),
    .A2(net541),
    .A3(net1072),
    .S0(net542),
    .S1(net532),
    .X(net543));
 sky130_fd_sc_hd__xnor2_1 c674 (.A(net540),
    .B(net425),
    .Y(net544));
 sky130_fd_sc_hd__buf_1 c675 (.A(net680),
    .X(net545));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net538),
    .A1(net541),
    .A2(net540),
    .A3(net431),
    .S0(net1023),
    .S1(net715),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_2 c677 (.A(net680),
    .X(net547));
 sky130_fd_sc_hd__xnor2_4 c678 (.A(net1014),
    .B(net877),
    .Y(net548));
 sky130_fd_sc_hd__xnor2_1 c679 (.A(net547),
    .B(net541),
    .Y(net549));
 sky130_fd_sc_hd__xnor2_2 c68 (.A(net4),
    .B(net917),
    .Y(net6));
 sky130_fd_sc_hd__a21bo_1 c680 (.A1(net549),
    .A2(net536),
    .B1_N(net540),
    .X(net550));
 sky130_fd_sc_hd__a41o_2 c681 (.A1(net549),
    .A2(net1014),
    .A3(net547),
    .A4(net715),
    .B1(net878),
    .X(net551));
 sky130_fd_sc_hd__a21bo_2 c682 (.A1(net196),
    .A2(net547),
    .B1_N(net447),
    .X(net552));
 sky130_fd_sc_hd__a31o_1 c683 (.A1(net445),
    .A2(net1014),
    .A3(net552),
    .B1(net1040),
    .X(net553));
 sky130_fd_sc_hd__a21bo_1 c684 (.A1(net550),
    .A2(net544),
    .B1_N(net547),
    .X(net554));
 sky130_fd_sc_hd__sdfrtp_4 c685 (.CLK(clknet_4_11_0_clk),
    .D(net1020),
    .RESET_B(net1078),
    .SCD(net554),
    .SCE(clknet_1_0__leaf_net866),
    .Q(net555));
 sky130_fd_sc_hd__mux4_2 c686 (.A0(net536),
    .A1(net1038),
    .A2(net544),
    .A3(net110),
    .S0(net1093),
    .S1(net865),
    .X(net556));
 sky130_fd_sc_hd__a31o_1 c687 (.A1(net541),
    .A2(net922),
    .A3(net550),
    .B1(net1012),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(net539),
    .A1(net551),
    .A2(net555),
    .A3(net536),
    .S0(net552),
    .S1(net865),
    .X(net558));
 sky130_fd_sc_hd__a31o_1 c689 (.A1(net1037),
    .A2(net1014),
    .A3(clknet_1_0__leaf_net846),
    .B1(net865),
    .X(net559));
 sky130_fd_sc_hd__xnor2_2 c69 (.A(net950),
    .B(net917),
    .Y(net7));
 sky130_fd_sc_hd__sdfbbp_1 c690 (.CLK(clknet_4_10_0_clk),
    .D(net537),
    .RESET_B(net1080),
    .SCD(net1012),
    .SCE(net533),
    .SET_B(net231),
    .Q(net561),
    .Q_N(net560));
 sky130_fd_sc_hd__sdfrtp_1 c691 (.CLK(clknet_4_10_0_clk),
    .D(net553),
    .RESET_B(net110),
    .SCD(net445),
    .SCE(net1012),
    .Q(net562));
 sky130_fd_sc_hd__a41o_2 c692 (.A1(net347),
    .A2(net547),
    .A3(net537),
    .A4(net1023),
    .B1(net551),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net554),
    .A1(net560),
    .A2(net552),
    .A3(net539),
    .S0(net1040),
    .S1(net865),
    .X(net564));
 sky130_fd_sc_hd__a31o_1 c694 (.A1(net237),
    .A2(net555),
    .A3(net561),
    .B1(net563),
    .X(net565));
 sky130_fd_sc_hd__sdfsbp_1 c695 (.CLK(clknet_4_11_0_clk),
    .D(net563),
    .SCD(net552),
    .SCE(net1012),
    .SET_B(net773),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__sdfbbn_1 c696 (.CLK_N(clknet_4_10_0_clk),
    .D(net562),
    .RESET_B(net539),
    .SCD(net237),
    .SCE(net445),
    .SET_B(clknet_1_1__leaf_net847),
    .Q(net569),
    .Q_N(net568));
 sky130_fd_sc_hd__sdfsbp_1 c697 (.CLK(clknet_4_11_0_clk),
    .D(net533),
    .SCD(net231),
    .SCE(net541),
    .SET_B(net1055),
    .Q(net571),
    .Q_N(net570));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(net1046),
    .A2(net562),
    .A3(net570),
    .B1(net554),
    .X(net572));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net569),
    .A1(net110),
    .A2(net541),
    .A3(net547),
    .S0(net567),
    .S1(net1038),
    .X(net573));
 sky130_fd_sc_hd__buf_4 c70 (.A(net709),
    .X(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net561),
    .A1(net430),
    .A2(net571),
    .A3(net569),
    .S0(net1012),
    .S1(net786),
    .X(net574));
 sky130_fd_sc_hd__a41o_1 c701 (.A1(net567),
    .A2(net562),
    .A3(net548),
    .A4(net774),
    .B1(net865),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net571),
    .A1(net575),
    .A2(net447),
    .A3(net1037),
    .S0(net774),
    .S1(net776),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net234),
    .A1(net575),
    .A2(net573),
    .A3(net1087),
    .S0(net568),
    .S1(net780),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net430),
    .A1(net231),
    .A2(net952),
    .A3(net552),
    .S0(net1012),
    .S1(net1032),
    .X(net578));
 sky130_fd_sc_hd__a41o_1 c705 (.A1(net448),
    .A2(net955),
    .A3(clknet_1_0__leaf_net477),
    .A4(net1014),
    .B1(net947),
    .X(net579));
 sky130_fd_sc_hd__a41o_1 c706 (.A1(net573),
    .A2(net1014),
    .A3(clknet_1_1__leaf_net579),
    .A4(net548),
    .B1(net1041),
    .X(net580));
 sky130_fd_sc_hd__sdfbbn_1 c707 (.CLK_N(clknet_4_11_0_clk),
    .D(net349),
    .RESET_B(net231),
    .SCD(clknet_1_0__leaf_net579),
    .SCE(net1012),
    .SET_B(net922),
    .Q(net582),
    .Q_N(net581));
 sky130_fd_sc_hd__a41o_1 c708 (.A1(net947),
    .A2(net582),
    .A3(net1012),
    .A4(clknet_1_1__leaf_net579),
    .B1(net881),
    .X(net583));
 sky130_fd_sc_hd__a41o_1 c709 (.A1(net1014),
    .A2(net904),
    .A3(net551),
    .A4(clknet_1_1__leaf_net579),
    .B1(net879),
    .X(net584));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net935),
    .B(net952),
    .Y(net9));
 sky130_fd_sc_hd__a41o_1 c710 (.A1(net342),
    .A2(net551),
    .A3(net430),
    .A4(clknet_1_0__leaf_net866),
    .B1(net880),
    .X(net585));
 sky130_fd_sc_hd__a41o_1 c711 (.A1(net575),
    .A2(net87),
    .A3(net551),
    .A4(net581),
    .B1(clknet_1_0__leaf_net579),
    .X(net586));
 sky130_fd_sc_hd__a41o_1 c712 (.A1(net582),
    .A2(net467),
    .A3(clknet_1_0__leaf_net579),
    .A4(clknet_1_0__leaf_net867),
    .B1(net880),
    .X(net587));
 sky130_fd_sc_hd__a41o_1 c713 (.A1(net559),
    .A2(clknet_1_1__leaf_net119),
    .A3(net551),
    .A4(net581),
    .B1(net1045),
    .X(net588));
 sky130_fd_sc_hd__a41o_1 c714 (.A1(clknet_1_1__leaf_net579),
    .A2(net587),
    .A3(net551),
    .A4(net89),
    .B1(net843),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net1012),
    .A1(net909),
    .A2(clknet_1_1__leaf_net579),
    .A3(net821),
    .S0(net1041),
    .S1(net881),
    .X(net590));
 sky130_fd_sc_hd__a41o_1 c716 (.A1(net584),
    .A2(clknet_1_0__leaf_net588),
    .A3(net573),
    .A4(net447),
    .B1(clknet_1_0__leaf_net867),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(clknet_1_1__leaf_net588),
    .A1(net947),
    .A2(net786),
    .A3(net821),
    .S0(clknet_1_0__leaf_net867),
    .S1(net1039),
    .X(net592));
 sky130_fd_sc_hd__a41o_1 c718 (.A1(net551),
    .A2(net1023),
    .A3(net1014),
    .A4(net1032),
    .B1(net786),
    .X(net593));
 sky130_fd_sc_hd__a41o_1 c719 (.A1(net1023),
    .A2(net575),
    .A3(clknet_1_1__leaf_net579),
    .A4(net818),
    .B1(net881),
    .X(net594));
 sky130_fd_sc_hd__xnor2_2 c72 (.A(net933),
    .B(net9),
    .Y(net10));
 sky130_fd_sc_hd__a41o_1 c720 (.A1(clknet_1_1__leaf_net588),
    .A2(net89),
    .A3(net781),
    .A4(net1041),
    .B1(net1039),
    .X(net595));
 sky130_fd_sc_hd__a41o_1 c721 (.A1(net901),
    .A2(net231),
    .A3(clknet_1_1__leaf_net966),
    .A4(net799),
    .B1(clknet_1_0__leaf_net867),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net593),
    .A1(clknet_1_0__leaf_net588),
    .A2(clknet_1_0__leaf_net585),
    .A3(net922),
    .S0(net947),
    .S1(clknet_1_0__leaf_net579),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net1045),
    .A1(net593),
    .A2(net773),
    .A3(net805),
    .S0(clknet_1_0__leaf_net867),
    .S1(net879),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net231),
    .A1(net467),
    .A2(net259),
    .A3(clknet_1_0__leaf_net579),
    .S0(net413),
    .S1(net805),
    .X(net599));
 sky130_fd_sc_hd__a41o_1 c725 (.A1(clknet_1_0__leaf_net579),
    .A2(net780),
    .A3(net800),
    .A4(net880),
    .B1(net883),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net548),
    .A1(net552),
    .A2(net800),
    .A3(net1041),
    .S0(clknet_1_1__leaf_net847),
    .S1(net1039),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net413),
    .A1(net1025),
    .A2(net485),
    .A3(net563),
    .S0(net782),
    .S1(net1039),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net563),
    .A1(net947),
    .A2(net448),
    .A3(net91),
    .S0(net1016),
    .S1(net873),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net477),
    .A1(net1023),
    .A2(net259),
    .A3(net1012),
    .S0(net808),
    .S1(net882),
    .X(net604));
 sky130_fd_sc_hd__xnor2_1 c73 (.A(net957),
    .B(net2),
    .Y(net11));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(clknet_1_1__leaf_net119),
    .A1(net413),
    .A2(net1023),
    .A3(net552),
    .S0(net849),
    .S1(net883),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(clknet_1_0__leaf_net119),
    .A1(net1025),
    .A2(net448),
    .A3(net1022),
    .S0(net490),
    .S1(net1016),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net563),
    .A1(net485),
    .A2(net1023),
    .A3(net552),
    .S0(net1090),
    .S1(net1054),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net556),
    .A1(net548),
    .A2(net1032),
    .A3(net799),
    .S0(net873),
    .S1(net882),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net552),
    .A1(net556),
    .A2(net264),
    .A3(net1022),
    .S0(net1032),
    .S1(net1039),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net264),
    .A1(net556),
    .A2(net1022),
    .A3(net1025),
    .S0(net1023),
    .S1(clknet_1_1__leaf_net866),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net1032),
    .A1(net1023),
    .A2(clknet_1_1__leaf_net605),
    .A3(net489),
    .S0(net817),
    .S1(net1039),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net1023),
    .A1(net1025),
    .A2(net307),
    .A3(net906),
    .S0(net796),
    .S1(net834),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net123),
    .A1(net612),
    .A2(net548),
    .A3(net898),
    .S0(clknet_1_1__leaf_net866),
    .S1(clknet_1_0__leaf_net885),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(clknet_1_1__leaf_net477),
    .A1(net1033),
    .A2(net563),
    .A3(net821),
    .S0(net1039),
    .S1(clknet_1_0__leaf_net885),
    .X(net614));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net2),
    .B(net9),
    .Y(net12));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net337),
    .A1(net1032),
    .A2(net1025),
    .A3(net819),
    .S0(net1039),
    .S1(clknet_1_0__leaf_net884),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net490),
    .A1(net548),
    .A2(net799),
    .A3(net1039),
    .S0(clknet_1_0__leaf_net884),
    .S1(clknet_1_0__leaf_net885),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_1__leaf_net616),
    .A1(net986),
    .A2(net786),
    .A3(net817),
    .S0(net1039),
    .S1(clknet_1_0__leaf_net885),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(clknet_1_0__leaf_net605),
    .A1(net545),
    .A2(net448),
    .A3(clknet_1_0__leaf_net616),
    .S0(net817),
    .S1(net833),
    .X(net618));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net123),
    .A1(net905),
    .A2(net739),
    .A3(net796),
    .S0(clknet_1_1__leaf_net884),
    .S1(clknet_1_0__leaf_net885),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net548),
    .A1(net1017),
    .A2(net781),
    .A3(net818),
    .S0(clknet_1_1__leaf_net885),
    .S1(clknet_1_1__leaf_net886),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net337),
    .A1(net413),
    .A2(clknet_1_1__leaf_net600),
    .A3(net806),
    .S0(net817),
    .S1(clknet_1_0__leaf_net886),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net601),
    .A1(net1037),
    .A2(net776),
    .A3(net806),
    .S0(clknet_1_0__leaf_net885),
    .S1(clknet_1_0__leaf_net886),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net1013),
    .A1(clknet_1_1__leaf_net409),
    .A2(clknet_1_1__leaf_net491),
    .A3(net943),
    .S0(clknet_1_0__leaf_net846),
    .S1(clknet_1_1__leaf_net885),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_0__leaf_net409),
    .A1(net555),
    .A2(net91),
    .A3(net1041),
    .S0(clknet_1_1__leaf_net885),
    .S1(net889),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 c75 (.A(net709),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net555),
    .A1(net89),
    .A2(net1013),
    .A3(clknet_1_1__leaf_net867),
    .S0(net873),
    .S1(net876),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net1026),
    .A1(net555),
    .A2(clknet_1_0__leaf_net409),
    .A3(net876),
    .S0(net888),
    .S1(net890),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(clknet_1_1__leaf_net491),
    .A1(net529),
    .A2(clknet_1_1__leaf_net409),
    .A3(net963),
    .S0(clknet_1_0__leaf_net846),
    .S1(net887),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(clknet_1_1__leaf_net585),
    .A1(clknet_1_0__leaf_net600),
    .A2(net529),
    .A3(net485),
    .S0(net922),
    .S1(net888),
    .X(net628));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net548),
    .A1(net361),
    .A2(clknet_1_1__leaf_net491),
    .A3(clknet_1_1__leaf_net409),
    .S0(net834),
    .S1(net891),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net490),
    .A1(clknet_1_1__leaf_net966),
    .A2(net1025),
    .A3(net819),
    .S0(clknet_1_0__leaf_net846),
    .S1(net892),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net361),
    .A1(clknet_1_1__leaf_net409),
    .A2(net487),
    .A3(net259),
    .S0(net922),
    .S1(net799),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net1025),
    .A1(net1013),
    .A2(clknet_1_1__leaf_net409),
    .A3(clknet_1_1__leaf_net867),
    .S0(net894),
    .S1(net895),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net580),
    .A1(net986),
    .A2(net91),
    .A3(net818),
    .S0(clknet_1_1__leaf_net885),
    .S1(net894),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net487),
    .A1(net171),
    .A2(net818),
    .A3(clknet_1_1__leaf_net867),
    .S0(net873),
    .S1(net894),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c76 (.A0(net917),
    .A1(net908),
    .A2(net949),
    .A3(net8),
    .S0(net12),
    .S1(net942),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net528),
    .A1(net808),
    .A2(net1041),
    .A3(clknet_1_0__leaf_net846),
    .S0(net893),
    .S1(net894),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net548),
    .A1(net1025),
    .A2(net1017),
    .A3(net808),
    .S0(net1068),
    .S1(net895),
    .X(net636));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net485),
    .A1(net635),
    .A2(net1025),
    .A3(net782),
    .S0(net801),
    .S1(net876),
    .X(net637));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net637),
    .A1(net1025),
    .A2(net123),
    .A3(net548),
    .S0(net802),
    .S1(net806),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net1017),
    .A1(net739),
    .A2(net801),
    .A3(net806),
    .S0(net876),
    .S1(net893),
    .X(net639));
 sky130_fd_sc_hd__xnor2_4 c77 (.A(net5),
    .B(net823),
    .Y(net15));
 sky130_fd_sc_hd__mux4_1 c78 (.A0(net945),
    .A1(net951),
    .A2(net954),
    .A3(net12),
    .S0(net15),
    .S1(net822),
    .X(net16));
 sky130_fd_sc_hd__xnor2_4 c79 (.A(net1043),
    .B(net8),
    .Y(net974));
 sky130_fd_sc_hd__xnor2_1 c80 (.A(net936),
    .B(net7),
    .Y(net17));
 sky130_fd_sc_hd__xnor2_1 c81 (.A(net17),
    .B(net810),
    .Y(net18));
 sky130_fd_sc_hd__mux4_1 c82 (.A0(net10),
    .A1(net7),
    .A2(net1043),
    .A3(net1021),
    .S0(net12),
    .S1(net15),
    .X(net19));
 sky130_fd_sc_hd__xnor2_1 c83 (.A(net17),
    .B(net942),
    .Y(net20));
 sky130_fd_sc_hd__clkbuf_1 c84 (.A(net709),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 c85 (.A0(net8),
    .A1(net1043),
    .A2(net21),
    .A3(net12),
    .S0(net915),
    .S1(net15),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c86 (.A0(net21),
    .A1(net11),
    .A2(net18),
    .A3(net13),
    .S0(net820),
    .S1(net824),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c87 (.A0(net940),
    .A1(net1043),
    .A2(net914),
    .A3(net1021),
    .S0(net825),
    .S1(net826),
    .X(net24));
 sky130_fd_sc_hd__xnor2_4 c88 (.A(net914),
    .B(net957),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_1 c89 (.A(net10),
    .B(net810),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net922),
    .B(net8),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_4 c91 (.A(net937),
    .B(net13),
    .Y(net28));
 sky130_fd_sc_hd__buf_1 c92 (.A(net714),
    .X(net29));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net951),
    .B(net27),
    .Y(net30));
 sky130_fd_sc_hd__sdfbbn_1 c94 (.CLK_N(clknet_4_4_0_clk),
    .D(net20),
    .RESET_B(net28),
    .SCD(net29),
    .SCE(net30),
    .SET_B(net824),
    .Q(net32),
    .Q_N(net31));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net30),
    .B(net1021),
    .Y(net33));
 sky130_fd_sc_hd__a21bo_1 c96 (.A1(net13),
    .A2(net27),
    .B1_N(net823),
    .X(net34));
 sky130_fd_sc_hd__a21bo_1 c97 (.A1(net29),
    .A2(net34),
    .B1_N(net30),
    .X(net35));
 sky130_fd_sc_hd__mux4_1 c98 (.A0(net35),
    .A1(net944),
    .A2(net34),
    .A3(net8),
    .S0(net33),
    .S1(net28),
    .X(net36));
 sky130_fd_sc_hd__a21bo_2 c99 (.A1(net32),
    .A2(net28),
    .B1_N(net1061),
    .X(net37));
 sky130_fd_sc_hd__a31o_1 merge765 (.A1(net207),
    .A2(net532),
    .A3(net208),
    .B1(net861),
    .X(net640));
 sky130_fd_sc_hd__a41o_1 merge766 (.A1(net246),
    .A2(net252),
    .A3(net75),
    .A4(clknet_1_0__leaf_net243),
    .B1(net231),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net916),
    .A1(clknet_1_0__leaf_net966),
    .A2(net18),
    .A3(net1036),
    .S0(net137),
    .S1(net829),
    .X(net642));
 sky130_fd_sc_hd__a31o_1 merge768 (.A1(clknet_1_1__leaf_net354),
    .A2(net330),
    .A3(net941),
    .B1(net850),
    .X(net643));
 sky130_fd_sc_hd__a31o_1 merge769 (.A1(net100),
    .A2(net75),
    .A3(net1),
    .B1(net124),
    .X(net644));
 sky130_fd_sc_hd__a41o_1 merge770 (.A1(net919),
    .A2(net74),
    .A3(net77),
    .A4(net73),
    .B1(net79),
    .X(net645));
 sky130_fd_sc_hd__mux4_1 merge771 (.A0(net96),
    .A1(net90),
    .A2(net95),
    .A3(net101),
    .S0(net941),
    .S1(net83),
    .X(net646));
 sky130_fd_sc_hd__a31o_1 merge772 (.A1(net1002),
    .A2(net52),
    .A3(net56),
    .B1(net1051),
    .X(net647));
 sky130_fd_sc_hd__a41o_1 merge773 (.A1(net27),
    .A2(net20),
    .A3(net42),
    .A4(net38),
    .B1(net1061),
    .X(net648));
 sky130_fd_sc_hd__a41o_1 merge774 (.A1(net330),
    .A2(net318),
    .A3(net85),
    .A4(net206),
    .B1(net1040),
    .X(net649));
 sky130_fd_sc_hd__a31o_1 merge775 (.A1(net166),
    .A2(net84),
    .A3(net168),
    .B1(net906),
    .X(net650));
 sky130_fd_sc_hd__a31o_1 merge776 (.A1(net144),
    .A2(net84),
    .A3(net6),
    .B1(net1076),
    .X(net651));
 sky130_fd_sc_hd__a31o_1 merge777 (.A1(net240),
    .A2(net340),
    .A3(clknet_1_0__leaf_net354),
    .B1(net848),
    .X(net652));
 sky130_fd_sc_hd__a31o_1 merge778 (.A1(net904),
    .A2(net207),
    .A3(net415),
    .B1(net414),
    .X(net653));
 sky130_fd_sc_hd__a41o_1 merge779 (.A1(net107),
    .A2(net1029),
    .A3(net907),
    .A4(net211),
    .B1(clknet_1_1__leaf_net828),
    .X(net654));
 sky130_fd_sc_hd__a31o_1 merge780 (.A1(net952),
    .A2(net84),
    .A3(net896),
    .B1(net90),
    .X(net655));
 sky130_fd_sc_hd__a31o_1 merge781 (.A1(net76),
    .A2(net218),
    .A3(net89),
    .B1(net1022),
    .X(net656));
 sky130_fd_sc_hd__a31o_1 merge782 (.A1(net6),
    .A2(net4),
    .A3(net11),
    .B1(net10),
    .X(net657));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(clknet_1_0__leaf_net966),
    .A1(net373),
    .A2(net982),
    .A3(net377),
    .S0(net794),
    .S1(net854),
    .X(net658));
 sky130_fd_sc_hd__a41o_1 merge784 (.A1(net439),
    .A2(net312),
    .A3(clknet_1_1__leaf_net845),
    .A4(clknet_1_0__leaf_net847),
    .B1(net863),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net73),
    .A1(net1000),
    .A2(net981),
    .A3(net182),
    .S0(net978),
    .S1(net835),
    .X(net660));
 sky130_fd_sc_hd__a31o_1 merge786 (.A1(clknet_1_1__leaf_net131),
    .A2(clknet_1_0__leaf_net353),
    .A3(clknet_1_1__leaf_net354),
    .B1(net831),
    .X(net661));
 sky130_fd_sc_hd__buf_1 merge787 (.A(clknet_1_0__leaf_net749),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_1 merge788 (.A(net815),
    .X(net663));
 sky130_fd_sc_hd__a31o_1 merge789 (.A1(net458),
    .A2(clknet_1_0__leaf_net354),
    .A3(net947),
    .B1(net352),
    .X(net664));
 sky130_fd_sc_hd__a41o_1 merge790 (.A1(net374),
    .A2(net377),
    .A3(net340),
    .A4(clknet_1_1__leaf_net380),
    .B1(net854),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net224),
    .A1(net283),
    .A2(net189),
    .A3(net141),
    .S0(net1034),
    .S1(net833),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net167),
    .A1(net163),
    .A2(net1013),
    .A3(net187),
    .S0(net25),
    .S1(net73),
    .X(net667));
 sky130_fd_sc_hd__a41o_1 merge793 (.A1(net4),
    .A2(net18),
    .A3(net104),
    .A4(net904),
    .B1(net100),
    .X(net668));
 sky130_fd_sc_hd__a41o_1 merge794 (.A1(clknet_1_1__leaf_net243),
    .A2(net256),
    .A3(net264),
    .A4(net248),
    .B1(net839),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_1 merge795 (.A(net816),
    .X(net670));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(clknet_1_1__leaf_net165),
    .A1(net992),
    .A2(net33),
    .A3(net1013),
    .S0(net710),
    .S1(net836),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 merge797 (.A0(clknet_1_1__leaf_net271),
    .A1(net123),
    .A2(net297),
    .A3(net960),
    .S0(net994),
    .S1(net820),
    .X(net672));
 sky130_fd_sc_hd__a41o_1 merge798 (.A1(net196),
    .A2(net84),
    .A3(net1057),
    .A4(net206),
    .B1(net90),
    .X(net673));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net211),
    .A1(net229),
    .A2(net224),
    .A3(net207),
    .S0(net200),
    .S1(net204),
    .X(net674));
 sky130_fd_sc_hd__a41o_1 merge800 (.A1(net439),
    .A2(net434),
    .A3(net437),
    .A4(net202),
    .B1(clknet_1_0__leaf_net847),
    .X(net675));
 sky130_fd_sc_hd__mux4_1 merge801 (.A0(net24),
    .A1(net139),
    .A2(net899),
    .A3(net168),
    .S0(net167),
    .S1(net705),
    .X(net676));
 sky130_fd_sc_hd__mux4_1 merge802 (.A0(net953),
    .A1(clknet_1_1__leaf_net243),
    .A2(net1019),
    .A3(clknet_1_1__leaf_net140),
    .S0(clknet_1_0__leaf_net966),
    .S1(net12),
    .X(net677));
 sky130_fd_sc_hd__mux4_1 merge803 (.A0(net74),
    .A1(net310),
    .A2(net1020),
    .A3(net914),
    .S0(net1081),
    .S1(net340),
    .X(net678));
 sky130_fd_sc_hd__mux4_1 merge804 (.A0(net324),
    .A1(net312),
    .A2(net457),
    .A3(net433),
    .S0(net348),
    .S1(net863),
    .X(net679));
 sky130_fd_sc_hd__sdfstp_1 merge805 (.CLK(clknet_4_10_0_clk),
    .D(net415),
    .SCD(net1022),
    .SCE(net431),
    .SET_B(net535),
    .Q(net680));
 sky130_fd_sc_hd__sdfbbp_1 merge806 (.CLK(clknet_4_8_0_clk),
    .D(net416),
    .RESET_B(net902),
    .SCD(net415),
    .SCE(net1033),
    .SET_B(net1056),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__mux4_1 merge807 (.A0(net242),
    .A1(net247),
    .A2(net246),
    .A3(net5),
    .S0(net144),
    .S1(net73),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 merge808 (.A0(net433),
    .A1(net250),
    .A2(net1015),
    .A3(net463),
    .S0(net434),
    .S1(net449),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 merge809 (.A0(net206),
    .A1(net996),
    .A2(net1029),
    .A3(clknet_1_0__leaf_net228),
    .S0(clknet_1_0__leaf_net233),
    .S1(net232),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 merge810 (.A0(net338),
    .A1(net333),
    .A2(net321),
    .A3(net322),
    .S0(net232),
    .S1(net1071),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 merge811 (.A0(net107),
    .A1(clknet_1_1__leaf_net228),
    .A2(net420),
    .A3(net434),
    .S0(net921),
    .S1(net743),
    .X(net687));
 sky130_fd_sc_hd__a41o_1 merge812 (.A1(net1002),
    .A2(net46),
    .A3(net45),
    .A4(net33),
    .B1(net824),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 merge813 (.A0(net139),
    .A1(clknet_1_0__leaf_net140),
    .A2(net954),
    .A3(net15),
    .S0(clknet_1_0__leaf_net142),
    .S1(net24),
    .X(net689));
 sky130_fd_sc_hd__mux4_1 merge814 (.A0(net444),
    .A1(net446),
    .A2(net434),
    .A3(net930),
    .S0(net74),
    .S1(net76),
    .X(net690));
 sky130_fd_sc_hd__mux4_1 merge815 (.A0(net423),
    .A1(net415),
    .A2(net317),
    .A3(net319),
    .S0(net315),
    .S1(net321),
    .X(net691));
 sky130_fd_sc_hd__mux4_1 merge816 (.A0(net915),
    .A1(net44),
    .A2(net56),
    .A3(net1045),
    .S0(net58),
    .S1(net810),
    .X(net692));
 sky130_fd_sc_hd__mux4_1 merge817 (.A0(net222),
    .A1(net215),
    .A2(net219),
    .A3(clknet_1_0__leaf_net358),
    .S0(clknet_1_0__leaf_net355),
    .S1(net1015),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 merge818 (.A0(net309),
    .A1(net208),
    .A2(net1029),
    .A3(net204),
    .S0(net222),
    .S1(net206),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 merge819 (.A0(net90),
    .A1(net1031),
    .A2(net34),
    .A3(net44),
    .S0(net39),
    .S1(net1084),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 merge820 (.A0(net209),
    .A1(clknet_1_1__leaf_net225),
    .A2(net110),
    .A3(clknet_1_1__leaf_net129),
    .S0(net255),
    .S1(net259),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 merge821 (.A0(net322),
    .A1(net319),
    .A2(net321),
    .A3(net218),
    .S0(net530),
    .S1(net200),
    .X(net697));
 sky130_fd_sc_hd__mux4_1 merge822 (.A0(net201),
    .A1(net312),
    .A2(net311),
    .A3(net535),
    .S0(net431),
    .S1(net1033),
    .X(net698));
 sky130_fd_sc_hd__sdfbbn_1 merge823 (.CLK_N(clknet_4_8_0_clk),
    .D(net418),
    .RESET_B(net1024),
    .SCD(net415),
    .SCE(net429),
    .SET_B(net1038),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dfrbp_1 merge824 (.CLK(clknet_4_5_0_clk),
    .D(net64),
    .RESET_B(net1052),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net372),
    .B(net382),
    .Y(net703));
 sky130_fd_sc_hd__dfrbp_1 merge826 (.CLK(clknet_4_1_0_clk),
    .D(net121),
    .RESET_B(net126),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net639),
    .B(net625),
    .Y(net706));
 sky130_fd_sc_hd__dfrtn_1 merge828 (.CLK_N(clknet_4_13_0_clk),
    .D(net507),
    .RESET_B(net508),
    .Q(net707));
 sky130_fd_sc_hd__dfrtp_1 merge829 (.CLK(clknet_4_0_0_clk),
    .D(net216),
    .RESET_B(net655),
    .Q(net708));
 sky130_fd_sc_hd__dfrtp_1 merge830 (.CLK(clknet_4_1_0_clk),
    .D(net657),
    .RESET_B(net668),
    .Q(net709));
 sky130_fd_sc_hd__dfrtp_2 merge831 (.CLK(clknet_4_5_0_clk),
    .D(net169),
    .RESET_B(net170),
    .Q(net710));
 sky130_fd_sc_hd__dfsbp_1 merge832 (.CLK(clknet_4_8_0_clk),
    .D(net426),
    .SET_B(net653),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__dfsbp_1 merge833 (.CLK(clknet_4_4_0_clk),
    .D(net648),
    .SET_B(net692),
    .Q(net714),
    .Q_N(net713));
 sky130_fd_sc_hd__dfstp_1 merge834 (.CLK(clknet_4_10_0_clk),
    .D(net531),
    .SET_B(net543),
    .Q(net715));
 sky130_fd_sc_hd__dfstp_1 merge835 (.CLK(clknet_4_9_0_clk),
    .D(net360),
    .SET_B(net368),
    .Q(net716));
 sky130_fd_sc_hd__dfstp_1 merge836 (.CLK(clknet_4_8_0_clk),
    .D(net656),
    .SET_B(net678),
    .Q(net717));
 sky130_fd_sc_hd__dlrbn_1 merge837 (.D(net649),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net686),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net558),
    .B(net565),
    .Y(net720));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net289),
    .B(net287),
    .Y(net721));
 sky130_fd_sc_hd__xnor2_1 merge840 (.A(net578),
    .B(net583),
    .Y(net722));
 sky130_fd_sc_hd__xnor2_1 merge841 (.A(net191),
    .B(net194),
    .Y(net723));
 sky130_fd_sc_hd__dlrbn_1 merge842 (.D(net268),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net269),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__xnor2_1 merge843 (.A(net149),
    .B(net154),
    .Y(net726));
 sky130_fd_sc_hd__xnor2_1 merge844 (.A(net480),
    .B(net497),
    .Y(net727));
 sky130_fd_sc_hd__xnor2_1 merge845 (.A(net226),
    .B(net241),
    .Y(net728));
 sky130_fd_sc_hd__xnor2_1 merge846 (.A(net257),
    .B(net263),
    .Y(net729));
 sky130_fd_sc_hd__xnor2_1 merge847 (.A(net459),
    .B(net470),
    .Y(net730));
 sky130_fd_sc_hd__dlrbp_1 merge848 (.D(net659),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net675),
    .Q(net732),
    .Q_N(net731));
 sky130_fd_sc_hd__dlrbp_1 merge849 (.D(net645),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net93),
    .Q(net734),
    .Q_N(net733));
 sky130_fd_sc_hd__xnor2_1 merge850 (.A(net112),
    .B(net114),
    .Y(net735));
 sky130_fd_sc_hd__xnor2_1 merge851 (.A(net391),
    .B(net397),
    .Y(net736));
 sky130_fd_sc_hd__xnor2_1 merge852 (.A(net602),
    .B(net603),
    .Y(net737));
 sky130_fd_sc_hd__dlrtn_1 merge853 (.GATE_N(clknet_4_5_0_clk),
    .RESET_B(net304),
    .Q(net305));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net156),
    .B(net157),
    .Y(net738));
 sky130_fd_sc_hd__dlrtn_1 merge855 (.D(net617),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net638),
    .Q(net739));
 sky130_fd_sc_hd__xnor2_1 merge856 (.A(net738),
    .B(net102),
    .Y(net740));
 sky130_fd_sc_hd__dlrtn_1 merge857 (.D(net676),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net667),
    .Q(net741));
 sky130_fd_sc_hd__dlrtp_1 merge858 (.D(net690),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net679),
    .Q(net742));
 sky130_fd_sc_hd__dlrtp_1 merge859 (.D(net113),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net646),
    .Q(net743));
 sky130_fd_sc_hd__dlrtp_1 merge860 (.D(net693),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net687),
    .Q(net744));
 sky130_fd_sc_hd__xnor2_1 merge861 (.A(net410),
    .B(net387),
    .Y(net745));
 sky130_fd_sc_hd__edfxbp_1 merge862 (.CLK(clknet_4_5_0_clk),
    .D(net723),
    .DE(net660),
    .Q(net1007),
    .Q_N(net746));
 sky130_fd_sc_hd__edfxtp_1 merge863 (.CLK(clknet_4_3_0_clk),
    .D(net383),
    .DE(net683),
    .Q(net747));
 sky130_fd_sc_hd__sdlclkp_1 merge864 (.CLK(clknet_4_1_0_clk),
    .GATE(net735),
    .SCE(net644),
    .GCLK(net748));
 sky130_fd_sc_hd__sdlclkp_2 merge865 (.CLK(clknet_4_12_0_clk),
    .GATE(net730),
    .SCE(net684),
    .GCLK(net749));
 sky130_fd_sc_hd__sdlclkp_4 merge866 (.CLK(clknet_4_5_0_clk),
    .GATE(net290),
    .SCE(net688),
    .GCLK(net750));
 sky130_fd_sc_hd__dfrbp_1 merge867 (.CLK(clknet_4_6_0_clk),
    .D(net294),
    .RESET_B(net284),
    .Q(net994),
    .Q_N(net751));
 sky130_fd_sc_hd__xnor2_1 merge868 (.A(net503),
    .B(net504),
    .Y(net752));
 sky130_fd_sc_hd__dfrbp_1 merge869 (.CLK(clknet_4_2_0_clk),
    .D(net729),
    .RESET_B(net1058),
    .Q(net754),
    .Q_N(net753));
 sky130_fd_sc_hd__dfrtn_1 merge870 (.CLK_N(clknet_4_2_0_clk),
    .D(net685),
    .RESET_B(net654),
    .Q(net755));
 sky130_fd_sc_hd__dfrtp_1 merge871 (.CLK(clknet_4_7_0_clk),
    .D(net518),
    .RESET_B(net400),
    .Q(net977));
 sky130_fd_sc_hd__dfrtp_1 merge872 (.CLK(clknet_4_7_0_clk),
    .D(net403),
    .RESET_B(net745),
    .Q(net993));
 sky130_fd_sc_hd__xnor2_1 merge873 (.A(net598),
    .B(net629),
    .Y(net756));
 sky130_fd_sc_hd__xnor2_1 merge874 (.A(net574),
    .B(net621),
    .Y(net757));
 sky130_fd_sc_hd__dfrtp_1 merge875 (.CLK(clknet_4_13_0_clk),
    .D(net524),
    .RESET_B(net512),
    .Q(net758));
 sky130_fd_sc_hd__dfsbp_1 merge876 (.CLK(clknet_4_7_0_clk),
    .D(net671),
    .SET_B(net736),
    .Q(net760),
    .Q_N(net759));
 sky130_fd_sc_hd__dfsbp_1 merge877 (.CLK(clknet_4_2_0_clk),
    .D(net728),
    .SET_B(net696),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__dfstp_1 merge878 (.CLK(clknet_4_4_0_clk),
    .D(net642),
    .SET_B(net689),
    .Q(net763));
 sky130_fd_sc_hd__xnor2_1 merge879 (.A(net604),
    .B(net628),
    .Y(net764));
 sky130_fd_sc_hd__xnor2_1 merge880 (.A(net596),
    .B(net576),
    .Y(net765));
 sky130_fd_sc_hd__xnor2_1 merge881 (.A(net591),
    .B(net618),
    .Y(net766));
 sky130_fd_sc_hd__xnor2_1 merge882 (.A(net595),
    .B(net594),
    .Y(net767));
 sky130_fd_sc_hd__xnor2_1 merge883 (.A(net526),
    .B(net521),
    .Y(net768));
 sky130_fd_sc_hd__dfstp_1 merge884 (.CLK(clknet_4_5_0_clk),
    .D(net173),
    .SET_B(net651),
    .Q(net769));
 sky130_fd_sc_hd__xnor2_1 merge885 (.A(net706),
    .B(net767),
    .Y(net770));
 sky130_fd_sc_hd__xnor2_1 merge886 (.A(net513),
    .B(net626),
    .Y(net771));
 sky130_fd_sc_hd__dfstp_1 merge887 (.CLK(clknet_4_13_0_clk),
    .D(net514),
    .SET_B(net520),
    .Q(net772));
 sky130_fd_sc_hd__dlrbn_1 merge888 (.D(net557),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net720),
    .Q(net774),
    .Q_N(net773));
 sky130_fd_sc_hd__dlrbn_1 merge889 (.D(net757),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net694),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__dlrbp_1 merge890 (.D(net726),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net695),
    .Q(net778),
    .Q_N(net777));
 sky130_fd_sc_hd__xnor2_1 merge891 (.A(net615),
    .B(net592),
    .Y(net779));
 sky130_fd_sc_hd__dlrbp_1 merge892 (.D(net766),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net765),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dlrtn_2 merge893 (.D(net640),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net756),
    .Q(net782));
 sky130_fd_sc_hd__dlrtn_1 merge894 (.D(net278),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net677),
    .Q(net783));
 sky130_fd_sc_hd__dlrtn_1 merge895 (.D(net674),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net672),
    .Q(net784));
 sky130_fd_sc_hd__dlrtp_2 merge896 (.D(net661),
    .GATE(clknet_4_12_0_clk),
    .RESET_B(net771),
    .Q(net963));
 sky130_fd_sc_hd__dlrtp_2 merge897 (.D(net277),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net666),
    .Q(net785));
 sky130_fd_sc_hd__dlrtp_1 merge898 (.D(net572),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net722),
    .Q(net786));
 sky130_fd_sc_hd__xnor2_1 merge899 (.A(net608),
    .B(net613),
    .Y(net787));
 sky130_fd_sc_hd__xnor2_1 merge900 (.A(net609),
    .B(net610),
    .Y(net788));
 sky130_fd_sc_hd__edfxbp_1 merge901 (.CLK(clknet_4_9_0_clk),
    .D(net691),
    .DE(net664),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__edfxtp_1 merge902 (.CLK(clknet_4_3_0_clk),
    .D(net384),
    .DE(net643),
    .Q(net791));
 sky130_fd_sc_hd__sdlclkp_1 merge903 (.CLK(clknet_4_9_0_clk),
    .GATE(net652),
    .SCE(net370),
    .GCLK(net792));
 sky130_fd_sc_hd__sdlclkp_2 merge904 (.CLK(clknet_4_7_0_clk),
    .GATE(net371),
    .SCE(net768),
    .GCLK(net793));
 sky130_fd_sc_hd__sdlclkp_4 merge905 (.CLK(clknet_4_7_0_clk),
    .GATE(net282),
    .SCE(net301),
    .GCLK(net984));
 sky130_fd_sc_hd__dfrbp_1 merge906 (.CLK(clknet_4_3_0_clk),
    .D(net641),
    .RESET_B(net703),
    .Q(net795),
    .Q_N(net794));
 sky130_fd_sc_hd__dfrbp_1 merge907 (.CLK(clknet_4_14_0_clk),
    .D(net658),
    .RESET_B(net787),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__dfrtn_1 merge908 (.CLK_N(clknet_4_6_0_clk),
    .D(net669),
    .RESET_B(net650),
    .Q(net798));
 sky130_fd_sc_hd__dfrtp_2 merge909 (.CLK(clknet_4_14_0_clk),
    .D(net770),
    .RESET_B(net607),
    .Q(net799));
 sky130_fd_sc_hd__dfrtp_4 merge910 (.CLK(clknet_4_14_0_clk),
    .D(net369),
    .RESET_B(net597),
    .Q(net800));
 sky130_fd_sc_hd__dfrtp_2 merge911 (.CLK(clknet_4_13_0_clk),
    .D(net493),
    .RESET_B(net636),
    .Q(net801));
 sky130_fd_sc_hd__dfsbp_1 merge912 (.CLK(clknet_4_12_0_clk),
    .D(net386),
    .SET_B(net752),
    .Q(net803),
    .Q_N(net802));
 sky130_fd_sc_hd__dfsbp_1 merge913 (.CLK(clknet_4_11_0_clk),
    .D(net586),
    .SET_B(net665),
    .Q(net805),
    .Q_N(net804));
 sky130_fd_sc_hd__dfstp_1 merge914 (.CLK(clknet_4_15_0_clk),
    .D(net620),
    .SET_B(net634),
    .Q(net806));
 sky130_fd_sc_hd__dfstp_4 merge915 (.CLK(clknet_4_0_0_clk),
    .D(net214),
    .SET_B(net740),
    .Q(net807));
 sky130_fd_sc_hd__dfstp_1 merge916 (.CLK(clknet_4_12_0_clk),
    .D(net498),
    .SET_B(net633),
    .Q(net808));
 sky130_fd_sc_hd__dlrbn_2 merge917 (.D(net16),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net192),
    .Q(net810),
    .Q_N(net809));
 sky130_fd_sc_hd__dlrbn_1 merge918 (.D(net136),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net133),
    .Q(net812),
    .Q_N(net811));
 sky130_fd_sc_hd__dlrbp_1 merge919 (.D(net375),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net393),
    .Q(net814),
    .Q_N(net813));
 sky130_fd_sc_hd__dlrbp_1 merge920 (.D(net698),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net697),
    .Q(net816),
    .Q_N(net815));
 sky130_fd_sc_hd__dlrtn_1 merge921 (.D(net614),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net788),
    .Q(net817));
 sky130_fd_sc_hd__dlrtn_1 merge922 (.D(net779),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net632),
    .Q(net818));
 sky130_fd_sc_hd__dlrtn_1 merge923 (.D(net727),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net764),
    .Q(net819));
 sky130_fd_sc_hd__dlrtp_2 merge924 (.D(net19),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net721),
    .Q(net820));
 sky130_fd_sc_hd__dlrtp_1 merge925 (.D(net589),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net737),
    .Q(net821));
 sky130_fd_sc_hd__dfxbp_2 s926 (.CLK(clknet_4_4_0_clk),
    .D(net14),
    .Q(net823),
    .Q_N(net822));
 sky130_fd_sc_hd__dfxbp_1 s927 (.CLK(clknet_4_4_0_clk),
    .D(net22),
    .Q(net825),
    .Q_N(net824));
 sky130_fd_sc_hd__dfxtp_1 s928 (.CLK(clknet_4_4_0_clk),
    .D(net23),
    .Q(net826));
 sky130_fd_sc_hd__dfxtp_1 s929 (.CLK(clknet_4_4_0_clk),
    .D(net36),
    .Q(net827));
 sky130_fd_sc_hd__dfxtp_2 s930 (.CLK(clknet_4_5_0_clk),
    .D(net41),
    .Q(net997));
 sky130_fd_sc_hd__dlclkp_1 s931 (.CLK(clknet_4_5_0_clk),
    .GATE(net48),
    .GCLK(net991));
 sky130_fd_sc_hd__dlclkp_2 s932 (.CLK(clknet_4_5_0_clk),
    .GATE(net65),
    .GCLK(net1006));
 sky130_fd_sc_hd__dlclkp_4 s933 (.CLK(clknet_4_1_0_clk),
    .GATE(net111),
    .GCLK(net828));
 sky130_fd_sc_hd__dlxbn_1 s934 (.D(net132),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net830),
    .Q_N(net829));
 sky130_fd_sc_hd__dlxbn_1 s935 (.D(net134),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net832),
    .Q_N(net831));
 sky130_fd_sc_hd__dlxbp_1 s936 (.D(net148),
    .GATE(clknet_4_4_0_clk),
    .Q(net834),
    .Q_N(net833));
 sky130_fd_sc_hd__dlxtn_2 s937 (.D(net152),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net835));
 sky130_fd_sc_hd__dlxtn_2 s938 (.D(net176),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net836));
 sky130_fd_sc_hd__dlxtn_1 s939 (.D(net217),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net837));
 sky130_fd_sc_hd__dlxtp_1 s940 (.D(net238),
    .GATE(clknet_4_2_0_clk),
    .Q(net838));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s941 (.D(net253),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net839));
 sky130_fd_sc_hd__dfxbp_1 s942 (.CLK(clknet_4_5_0_clk),
    .D(net302),
    .Q(net964),
    .Q_N(net840));
 sky130_fd_sc_hd__dfxbp_1 s943 (.CLK(clknet_4_7_0_clk),
    .D(net303),
    .Q(net1003),
    .Q_N(net841));
 sky130_fd_sc_hd__dfxtp_1 s944 (.CLK(clknet_4_8_0_clk),
    .D(net325),
    .Q(net842));
 sky130_fd_sc_hd__dfxtp_1 s945 (.CLK(clknet_4_8_0_clk),
    .D(net326),
    .Q(net843));
 sky130_fd_sc_hd__dfxtp_1 s946 (.CLK(clknet_4_8_0_clk),
    .D(net336),
    .Q(net844));
 sky130_fd_sc_hd__dlclkp_1 s947 (.CLK(clknet_4_9_0_clk),
    .GATE(net339),
    .GCLK(net845));
 sky130_fd_sc_hd__dlclkp_2 s948 (.CLK(clknet_4_9_0_clk),
    .GATE(net341),
    .GCLK(net846));
 sky130_fd_sc_hd__dlclkp_4 s949 (.CLK(clknet_4_9_0_clk),
    .GATE(net344),
    .GCLK(net847));
 sky130_fd_sc_hd__dlxbn_1 s950 (.D(net346),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net849),
    .Q_N(net848));
 sky130_fd_sc_hd__dlxbn_1 s951 (.D(net362),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net851),
    .Q_N(net850));
 sky130_fd_sc_hd__dlxbp_1 s952 (.D(net364),
    .GATE(clknet_4_9_0_clk),
    .Q(net853),
    .Q_N(net852));
 sky130_fd_sc_hd__dlxtn_2 s953 (.D(net365),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net854));
 sky130_fd_sc_hd__dlxtn_1 s954 (.D(net388),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net855));
 sky130_fd_sc_hd__dlxtn_1 s955 (.D(net399),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net856));
 sky130_fd_sc_hd__dlxtp_1 s956 (.D(net406),
    .GATE(clknet_4_7_0_clk),
    .Q(net857));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s957 (.D(net411),
    .SLEEP_B(clknet_4_7_0_clk),
    .Q(net858));
 sky130_fd_sc_hd__dfxbp_1 s958 (.CLK(clknet_4_8_0_clk),
    .D(net419),
    .Q(net860),
    .Q_N(net859));
 sky130_fd_sc_hd__dfxbp_1 s959 (.CLK(clknet_4_8_0_clk),
    .D(net422),
    .Q(net862),
    .Q_N(net861));
 sky130_fd_sc_hd__dfxtp_1 s960 (.CLK(clknet_4_10_0_clk),
    .D(net442),
    .Q(net863));
 sky130_fd_sc_hd__dfxtp_1 s961 (.CLK(clknet_4_9_0_clk),
    .D(net450),
    .Q(net864));
 sky130_fd_sc_hd__dfxtp_1 s962 (.CLK(clknet_4_11_0_clk),
    .D(net454),
    .Q(net865));
 sky130_fd_sc_hd__dlclkp_1 s963 (.CLK(clknet_4_11_0_clk),
    .GATE(net456),
    .GCLK(net866));
 sky130_fd_sc_hd__dlclkp_2 s964 (.CLK(clknet_4_14_0_clk),
    .GATE(net472),
    .GCLK(net867));
 sky130_fd_sc_hd__dlclkp_4 s965 (.CLK(clknet_4_12_0_clk),
    .GATE(net474),
    .GCLK(net961));
 sky130_fd_sc_hd__dlxbn_1 s966 (.D(net475),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net869),
    .Q_N(net868));
 sky130_fd_sc_hd__dlxbn_2 s967 (.D(net494),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net990),
    .Q_N(net870));
 sky130_fd_sc_hd__dlxbp_1 s968 (.D(net495),
    .GATE(clknet_4_14_0_clk),
    .Q(net872),
    .Q_N(net871));
 sky130_fd_sc_hd__dlxtn_2 s969 (.D(net502),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net873));
 sky130_fd_sc_hd__dlxtn_4 s970 (.D(net516),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net980));
 sky130_fd_sc_hd__dlxtn_1 s971 (.D(net517),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net874));
 sky130_fd_sc_hd__dlxtp_1 s972 (.D(net522),
    .GATE(clknet_4_7_0_clk),
    .Q(net875));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s973 (.D(net527),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dfxbp_1 s974 (.CLK(clknet_4_10_0_clk),
    .D(net546),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dfxbp_1 s975 (.CLK(clknet_4_11_0_clk),
    .D(net564),
    .Q(net880),
    .Q_N(net879));
 sky130_fd_sc_hd__dfxtp_1 s976 (.CLK(clknet_4_11_0_clk),
    .D(net577),
    .Q(net881));
 sky130_fd_sc_hd__dfxtp_1 s977 (.CLK(clknet_4_14_0_clk),
    .D(net590),
    .Q(net882));
 sky130_fd_sc_hd__dfxtp_1 s978 (.CLK(clknet_4_14_0_clk),
    .D(net599),
    .Q(net883));
 sky130_fd_sc_hd__dlclkp_1 s979 (.CLK(clknet_4_14_0_clk),
    .GATE(net606),
    .GCLK(net884));
 sky130_fd_sc_hd__dlclkp_2 s980 (.CLK(clknet_4_14_0_clk),
    .GATE(net611),
    .GCLK(net885));
 sky130_fd_sc_hd__dlclkp_4 s981 (.CLK(clknet_4_15_0_clk),
    .GATE(net619),
    .GCLK(net886));
 sky130_fd_sc_hd__dlxbn_1 s982 (.D(net622),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__dlxbn_1 s983 (.D(net623),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net890),
    .Q_N(net889));
 sky130_fd_sc_hd__dlxbp_1 s984 (.D(net624),
    .GATE(clknet_4_15_0_clk),
    .Q(net892),
    .Q_N(net891));
 sky130_fd_sc_hd__dlxtn_1 s985 (.D(net627),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net893));
 sky130_fd_sc_hd__dlxtn_1 s986 (.D(net630),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net894));
 sky130_fd_sc_hd__dlxtn_1 s987 (.D(net631),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net895));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(in10),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in14),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net904));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net907));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net908));
 sky130_fd_sc_hd__buf_4 input14 (.A(in20),
    .X(net909));
 sky130_fd_sc_hd__buf_4 input15 (.A(in21),
    .X(net910));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net911));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in24),
    .X(net913));
 sky130_fd_sc_hd__buf_4 input19 (.A(in25),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net917));
 sky130_fd_sc_hd__buf_2 input23 (.A(in29),
    .X(net918));
 sky130_fd_sc_hd__buf_1 input24 (.A(in3),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net920));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_8 input27 (.A(in32),
    .X(net922));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(in33),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net924));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in36),
    .X(net926));
 sky130_fd_sc_hd__buf_2 input32 (.A(in37),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(in38),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in39),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net930));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net931));
 sky130_fd_sc_hd__buf_1 input37 (.A(in41),
    .X(net932));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net933));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(in43),
    .X(net934));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net935));
 sky130_fd_sc_hd__buf_1 input41 (.A(in45),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in46),
    .X(net937));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net938));
 sky130_fd_sc_hd__dlymetal6s2s_1 input44 (.A(in48),
    .X(net939));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in5),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(in50),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net943));
 sky130_fd_sc_hd__buf_1 input49 (.A(in52),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net945));
 sky130_fd_sc_hd__buf_1 input51 (.A(in54),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(in55),
    .X(net947));
 sky130_fd_sc_hd__buf_1 input53 (.A(in56),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(in57),
    .X(net949));
 sky130_fd_sc_hd__buf_1 input55 (.A(in58),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in59),
    .X(net951));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net952));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net954));
 sky130_fd_sc_hd__buf_4 input60 (.A(in7),
    .X(net955));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(in8),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(in9),
    .X(net957));
 sky130_fd_sc_hd__buf_2 output63 (.A(net958),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net959),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output65 (.A(net960),
    .X(out10));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(clknet_1_1__leaf_net961),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output67 (.A(net962),
    .X(out12));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net963),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output69 (.A(net964),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(clknet_1_0__leaf_net965),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(clknet_1_0__leaf_net966),
    .X(out16));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net967),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output73 (.A(net968),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net969),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output75 (.A(net970),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(clknet_1_1__leaf_net971),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output77 (.A(net972),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(clknet_1_1__leaf_net973),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output79 (.A(net1021),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output80 (.A(net975),
    .X(out24));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net976),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output82 (.A(net977),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output83 (.A(net978),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output84 (.A(net1018),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output85 (.A(net980),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output86 (.A(net981),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output87 (.A(net982),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output88 (.A(net983),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(clknet_1_1__leaf_net984),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output90 (.A(net985),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net986),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output92 (.A(net987),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output93 (.A(net988),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output94 (.A(net989),
    .X(out39));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net990),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(clknet_1_1__leaf_net991),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net992),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output98 (.A(net993),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net994),
    .X(out43));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(clknet_1_1__leaf_net995),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net996),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output102 (.A(net997),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output103 (.A(net998),
    .X(out49));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net999),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output105 (.A(net1000),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(clknet_1_1__leaf_net1001),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output107 (.A(net1002),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output108 (.A(net1003),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output109 (.A(net1004),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output110 (.A(net1005),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(clknet_1_0__leaf_net1006),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output112 (.A(net1007),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output113 (.A(net1008),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output114 (.A(net1034),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net1010),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output116 (.A(net1011),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net556),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net171),
    .X(net1013));
 sky130_fd_sc_hd__buf_4 max_cap119 (.A(net542),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net361),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net361),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net979),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 max_cap124 (.A(net958),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net202),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net974),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net307),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net545),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net424),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net967),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net967),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net970),
    .X(net1027));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net1031),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net198),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net198),
    .X(net1033));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net1009),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net98),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net87),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_4 fanout144 (.A(net882),
    .X(net1039));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net843),
    .X(net1040));
 sky130_fd_sc_hd__buf_4 max_cap146 (.A(net839),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_4 max_cap147 (.A(net838),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 max_cap148 (.A(net9),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 max_cap149 (.A(net92),
    .X(net1044));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net943),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net886 (.A(net886),
    .X(clknet_0_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_0__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net886 (.A(clknet_0_net886),
    .X(clknet_1_1__leaf_net886));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net885 (.A(net885),
    .X(clknet_0_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_0__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_1__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net961 (.A(net961),
    .X(clknet_0_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net477 (.A(net477),
    .X(clknet_0_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_0__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net477 (.A(clknet_0_net477),
    .X(clknet_1_1__leaf_net477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net579 (.A(net579),
    .X(clknet_0_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_0__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_1__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net476 (.A(net476),
    .X(clknet_0_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net491 (.A(net491),
    .X(clknet_0_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_0__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net491 (.A(clknet_0_net491),
    .X(clknet_1_1__leaf_net491));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net867 (.A(net867),
    .X(clknet_0_net867));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net867 (.A(clknet_0_net867),
    .X(clknet_1_0__leaf_net867));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net867 (.A(clknet_0_net867),
    .X(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net500 (.A(net500),
    .X(clknet_0_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_0__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_1__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net866 (.A(net866),
    .X(clknet_0_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_0__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net866 (.A(clknet_0_net866),
    .X(clknet_1_1__leaf_net866));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net847 (.A(net847),
    .X(clknet_0_net847));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net847 (.A(clknet_0_net847),
    .X(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net847 (.A(clknet_0_net847),
    .X(clknet_1_1__leaf_net847));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net358 (.A(net358),
    .X(clknet_0_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_0__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net358 (.A(clknet_0_net358),
    .X(clknet_1_1__leaf_net358));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net792 (.A(net792),
    .X(clknet_0_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net792 (.A(clknet_0_net792),
    .X(clknet_1_0__leaf_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net792 (.A(clknet_0_net792),
    .X(clknet_1_1__leaf_net792));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net355 (.A(net355),
    .X(clknet_0_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_0__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net355 (.A(clknet_0_net355),
    .X(clknet_1_1__leaf_net355));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net350 (.A(net350),
    .X(clknet_0_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_0__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net350 (.A(clknet_0_net350),
    .X(clknet_1_1__leaf_net350));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net353 (.A(net353),
    .X(clknet_0_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_0__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net353 (.A(clknet_0_net353),
    .X(clknet_1_1__leaf_net353));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net354 (.A(net354),
    .X(clknet_0_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_0__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net354 (.A(clknet_0_net354),
    .X(clknet_1_1__leaf_net354));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net846 (.A(net846),
    .X(clknet_0_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net846 (.A(clknet_0_net846),
    .X(clknet_1_1__leaf_net846));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net588 (.A(net588),
    .X(clknet_0_net588));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net588 (.A(clknet_0_net588),
    .X(clknet_1_0__leaf_net588));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net588 (.A(clknet_0_net588),
    .X(clknet_1_1__leaf_net588));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net845 (.A(net845),
    .X(clknet_0_net845));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net845 (.A(clknet_0_net845),
    .X(clknet_1_0__leaf_net845));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net845 (.A(clknet_0_net845),
    .X(clknet_1_1__leaf_net845));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net451 (.A(net451),
    .X(clknet_0_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_0__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net451 (.A(clknet_0_net451),
    .X(clknet_1_1__leaf_net451));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net455 (.A(net455),
    .X(clknet_0_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net828 (.A(net828),
    .X(clknet_0_net828));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net828 (.A(clknet_0_net828),
    .X(clknet_1_0__leaf_net828));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net828 (.A(clknet_0_net828),
    .X(clknet_1_1__leaf_net828));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net223 (.A(net223),
    .X(clknet_0_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_0__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net223 (.A(clknet_0_net223),
    .X(clknet_1_1__leaf_net223));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net254 (.A(net254),
    .X(clknet_0_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_1__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net228 (.A(net228),
    .X(clknet_0_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_0__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net228 (.A(clknet_0_net228),
    .X(clknet_1_1__leaf_net228));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net225 (.A(net225),
    .X(clknet_0_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_0__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_1__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net748 (.A(net748),
    .X(clknet_0_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net748 (.A(clknet_0_net748),
    .X(clknet_1_0__leaf_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net748 (.A(clknet_0_net748),
    .X(clknet_1_1__leaf_net748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net130 (.A(net130),
    .X(clknet_0_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_0__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net130 (.A(clknet_0_net130),
    .X(clknet_1_1__leaf_net130));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net125 (.A(net125),
    .X(clknet_0_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_0__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net125 (.A(clknet_0_net125),
    .X(clknet_1_1__leaf_net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net271 (.A(net271),
    .X(clknet_0_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net271 (.A(clknet_0_net271),
    .X(clknet_1_0__leaf_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net271 (.A(clknet_0_net271),
    .X(clknet_1_1__leaf_net271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net243 (.A(net243),
    .X(clknet_0_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_0__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_1__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net118 (.A(net118),
    .X(clknet_0_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_0__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net118 (.A(clknet_0_net118),
    .X(clknet_1_1__leaf_net118));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net131 (.A(net131),
    .X(clknet_0_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_0__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_1__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net127 (.A(net127),
    .X(clknet_0_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_0__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net127 (.A(clknet_0_net127),
    .X(clknet_1_1__leaf_net127));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net119 (.A(net119),
    .X(clknet_0_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net119 (.A(clknet_0_net119),
    .X(clknet_1_1__leaf_net119));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net143 (.A(net143),
    .X(clknet_0_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_0__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net143 (.A(clknet_0_net143),
    .X(clknet_1_1__leaf_net143));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net984 (.A(net984),
    .X(clknet_0_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_0__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net984 (.A(clknet_0_net984),
    .X(clknet_1_1__leaf_net984));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net404 (.A(net404),
    .X(clknet_0_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_0__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net404 (.A(clknet_0_net404),
    .X(clknet_1_1__leaf_net404));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net793 (.A(net793),
    .X(clknet_0_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_0__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net793 (.A(clknet_0_net793),
    .X(clknet_1_1__leaf_net793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net971 (.A(net971),
    .X(clknet_0_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_0__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net971 (.A(clknet_0_net971),
    .X(clknet_1_1__leaf_net971));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net389 (.A(net389),
    .X(clknet_0_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_0__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net389 (.A(clknet_0_net389),
    .X(clknet_1_1__leaf_net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net381 (.A(net381),
    .X(clknet_0_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_0__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net381 (.A(clknet_0_net381),
    .X(clknet_1_1__leaf_net381));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net379 (.A(net379),
    .X(clknet_0_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_0__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net379 (.A(clknet_0_net379),
    .X(clknet_1_1__leaf_net379));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net407 (.A(net407),
    .X(clknet_0_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_0__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net407 (.A(clknet_0_net407),
    .X(clknet_1_1__leaf_net407));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net966 (.A(net966),
    .X(clknet_0_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net966 (.A(clknet_0_net966),
    .X(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1006 (.A(net1006),
    .X(clknet_0_net1006));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1006 (.A(clknet_0_net1006),
    .X(clknet_1_0__leaf_net1006));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1006 (.A(clknet_0_net1006),
    .X(clknet_1_1__leaf_net1006));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net995 (.A(net995),
    .X(clknet_0_net995));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net995 (.A(clknet_0_net995),
    .X(clknet_1_0__leaf_net995));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net995 (.A(clknet_0_net995),
    .X(clknet_1_1__leaf_net995));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net965 (.A(net965),
    .X(clknet_0_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_0__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net965 (.A(clknet_0_net965),
    .X(clknet_1_1__leaf_net965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net991 (.A(net991),
    .X(clknet_0_net991));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net991 (.A(clknet_0_net991),
    .X(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net991 (.A(clknet_0_net991),
    .X(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net1001 (.A(net1001),
    .X(clknet_0_net1001));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net1001 (.A(clknet_0_net1001),
    .X(clknet_1_0__leaf_net1001));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net1001 (.A(clknet_0_net1001),
    .X(clknet_1_1__leaf_net1001));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net973 (.A(net973),
    .X(clknet_0_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net973 (.A(clknet_0_net973),
    .X(clknet_1_0__leaf_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net973 (.A(clknet_0_net973),
    .X(clknet_1_1__leaf_net973));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net164 (.A(net164),
    .X(clknet_0_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_1__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net750 (.A(net750),
    .X(clknet_0_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_0__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net750 (.A(clknet_0_net750),
    .X(clknet_1_1__leaf_net750));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net51 (.A(net51),
    .X(clknet_0_net51));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net51 (.A(clknet_0_net51),
    .X(clknet_1_0__leaf_net51));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net51 (.A(clknet_0_net51),
    .X(clknet_1_1__leaf_net51));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net47 (.A(net47),
    .X(clknet_0_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net47 (.A(clknet_0_net47),
    .X(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net47 (.A(clknet_0_net47),
    .X(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net749 (.A(net749),
    .X(clknet_0_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net749 (.A(clknet_0_net749),
    .X(clknet_1_0__leaf_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net749 (.A(clknet_0_net749),
    .X(clknet_1_1__leaf_net749));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net662 (.A(net662),
    .X(clknet_0_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_0__leaf_net662));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net662 (.A(clknet_0_net662),
    .X(clknet_1_1__leaf_net662));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net425),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net425),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net775),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net264),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net857),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net824),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net647),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net215),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net872),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net879),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net859),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net77),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net673),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net120),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net822),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net827),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net823),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net743),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net1042),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net855),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net835),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net852),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net876),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net854),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net715),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net844),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net536),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net836),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net731),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net841),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net39),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net81),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net552),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net60),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net555),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net236),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net758),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net702),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net829),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net833),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net874),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net566),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net861),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net424),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net821),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net840),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net363),
    .X(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_Q (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_Y (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_Y (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_SCE (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A4 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1_N (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S0 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_D (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1_N (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A4 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Y (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold8_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_RESET_B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_Q (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A4 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A3 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_RESET_B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_SCD (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SET_B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SET_B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_S1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_D (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCE (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_SCD (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_Q (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_S1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A3 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCE (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q_N (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_Q (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_RESET_B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_Q_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCD (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_Q (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_B1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A4 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_Q_N (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_S1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_Y (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A3 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_SCD (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_Q (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_Y (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_A4 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_Y (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_X (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_S1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_RESET_B (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A4 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_X (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_S0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_Q_N (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_D (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_Q (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_Y (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_Q (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SCD (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_Y (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_X (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_Y (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_A3 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_X (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_SCE (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Y (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_RESET_B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_Q (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_Q (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_Q (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A4 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_X (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_Q_N (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_Q (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A4 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_Y (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCD (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_X (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_Q (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_D (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_B1 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_X (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_Y (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_SET_B (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_D (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_D (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_Y (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_S1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A4 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_SCE (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_SCE (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_RESET_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_RESET_B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_D (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_SCE (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_A3 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_SCE (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_SCD (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_Y (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_B1_N (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_B1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_S1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A4 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_SCD (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_Q (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_Q_N (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_Q (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_S0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_Q (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge897_Q (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_RESET_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_Y (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_Q (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCD (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_Q (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A4 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge910_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A4 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_Q (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_Q_N (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_Q (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_SCE (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1_N (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge916_Q (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_Q (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge918_Q_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1_N (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge918_Q (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCE (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCD (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge923_Q (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A4 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge924_Q (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_B1_N (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_B1_N (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_Q (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B1_N (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_B1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_SCE (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B1_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A4 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCE (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCE (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_Q (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B1_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1_N (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_B1_N (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_B1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap146_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_s941_Q (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_SCE (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_D (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_B1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_Q (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net846_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_GCLK (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_Q (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A4 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_s969_Q (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A4 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A4 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_SCD (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_Q_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_Q (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_SCD (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A4 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A4 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_B1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B1_N (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A3 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_B1_N (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_SCE (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SET_B (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCD (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_SCD (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_D (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_A3 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_D (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_RESET_B (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_B1_N (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_D (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_RESET_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_Y (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCE (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_Q (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net966_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_DE (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_Q (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SCD (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_Q (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_Y (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_DE (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_A2 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_s970_Q (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A4 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_B1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCD (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SCE (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_DE (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_Q (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_B1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_SCD (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B1_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_Q (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_Q (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_S0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_B1_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_B1_N (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_S1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_RESET_B (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_SCD (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_SCE (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_SCE (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCE (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_SCD (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap119_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A4 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SCE (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_SCD (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_SCD (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_SCE (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1_N (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_D (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCD (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_D (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCD (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B1_N (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_SCD (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A4 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_RESET_B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_RESET_B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_RESET_B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SET_B (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCD (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A4 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SET_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_S1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_SCE (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_B1_N (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1_N (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCD (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B1_N (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_S1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B1_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1_N (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_B1_N (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_S1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_SET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_SET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_B1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_SCE (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_SCD (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_B1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_B1_N (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap146_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A4 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap147_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_SET_B (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_SCE (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_X (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_SCD (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_A3 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1_N (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge918_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge924_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge908_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge919_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge897_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge905_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_SLEEP_B (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s972_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge901_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge903_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge892_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge925_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s962_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s963_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s975_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s976_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_GATE (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge916_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s965_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s966_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s967_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge910_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge921_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s964_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s968_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s977_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s978_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s979_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s980_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge922_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s981_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s982_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s983_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s984_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s985_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s986_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s987_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net867_X (.DIODE(clknet_1_1__leaf_net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A4 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_B1 (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net847_X (.DIODE(clknet_1_0__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_S1 (.DIODE(clknet_1_1__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_SET_B (.DIODE(clknet_1_1__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(clknet_1_1__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net847_X (.DIODE(clknet_1_1__leaf_net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_B1 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A3 (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net846_X (.DIODE(clknet_1_0__leaf_net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net409_X (.DIODE(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net119_X (.DIODE(clknet_1_0__leaf_net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net966_A (.DIODE(clknet_0_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net966_A (.DIODE(clknet_0_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net966_X (.DIODE(clknet_0_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A1 (.DIODE(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A0 (.DIODE(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_S0 (.DIODE(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net966_X (.DIODE(clknet_1_0__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A0 (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_SCE (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net966_X (.DIODE(clknet_1_1__leaf_net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S1 (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1 (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net991_X (.DIODE(clknet_1_0__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_B (.DIODE(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_B1_N (.DIODE(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net991_X (.DIODE(clknet_1_1__leaf_net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_S1 (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_SCD (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_RESET_B (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net164_X (.DIODE(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_SET_B (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_D (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold8_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net212));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net425),
    .X(net1093));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
