module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net618;
 wire net671;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net798;
 wire clknet_1_0__leaf_net798;
 wire clknet_1_1__leaf_net798;
 wire clknet_0_net797;
 wire clknet_1_0__leaf_net797;
 wire clknet_1_1__leaf_net797;
 wire clknet_0_net796;
 wire clknet_1_0__leaf_net796;
 wire clknet_1_1__leaf_net796;
 wire clknet_0_net591;
 wire clknet_1_0__leaf_net591;
 wire clknet_1_1__leaf_net591;
 wire clknet_0_net565;
 wire clknet_1_0__leaf_net565;
 wire clknet_1_1__leaf_net565;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net779;
 wire clknet_1_0__leaf_net779;
 wire clknet_1_1__leaf_net779;
 wire clknet_0_net778;
 wire clknet_1_0__leaf_net778;
 wire clknet_1_1__leaf_net778;
 wire clknet_0_net777;
 wire clknet_1_0__leaf_net777;
 wire clknet_1_1__leaf_net777;
 wire clknet_0_net760;
 wire clknet_1_0__leaf_net760;
 wire clknet_1_1__leaf_net760;
 wire clknet_0_net479;
 wire clknet_1_0__leaf_net479;
 wire clknet_1_1__leaf_net479;
 wire clknet_0_net457;
 wire clknet_1_0__leaf_net457;
 wire clknet_1_1__leaf_net457;
 wire clknet_0_net458;
 wire clknet_1_0__leaf_net458;
 wire clknet_1_1__leaf_net458;
 wire clknet_0_net435;
 wire clknet_1_0__leaf_net435;
 wire clknet_1_1__leaf_net435;
 wire clknet_0_net546;
 wire clknet_1_0__leaf_net546;
 wire clknet_1_1__leaf_net546;
 wire clknet_0_net538;
 wire clknet_1_0__leaf_net538;
 wire clknet_1_1__leaf_net538;
 wire clknet_0_net703;
 wire clknet_1_0__leaf_net703;
 wire clknet_1_1__leaf_net703;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net471;
 wire clknet_1_0__leaf_net471;
 wire clknet_1_1__leaf_net471;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net542;
 wire clknet_1_0__leaf_net542;
 wire clknet_1_1__leaf_net542;
 wire clknet_0_net557;
 wire clknet_1_0__leaf_net557;
 wire clknet_1_1__leaf_net557;
 wire clknet_0_net559;
 wire clknet_1_0__leaf_net559;
 wire clknet_1_1__leaf_net559;
 wire clknet_0_net554;
 wire clknet_1_0__leaf_net554;
 wire clknet_1_1__leaf_net554;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net889;
 wire clknet_1_0__leaf_net889;
 wire clknet_1_1__leaf_net889;
 wire clknet_0_net378;
 wire clknet_1_0__leaf_net378;
 wire clknet_1_1__leaf_net378;
 wire clknet_0_net906;
 wire clknet_1_0__leaf_net906;
 wire clknet_1_1__leaf_net906;
 wire clknet_0_net919;
 wire clknet_1_0__leaf_net919;
 wire clknet_1_1__leaf_net919;
 wire clknet_0_net891;
 wire clknet_1_0__leaf_net891;
 wire clknet_1_1__leaf_net891;
 wire clknet_0_net743;
 wire clknet_1_0__leaf_net743;
 wire clknet_1_1__leaf_net743;
 wire clknet_0_net162;
 wire clknet_1_0__leaf_net162;
 wire clknet_1_1__leaf_net162;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net742;
 wire clknet_1_0__leaf_net742;
 wire clknet_1_1__leaf_net742;
 wire clknet_0_net256;
 wire clknet_1_0__leaf_net256;
 wire clknet_1_1__leaf_net256;
 wire clknet_0_net283;
 wire clknet_1_0__leaf_net283;
 wire clknet_1_1__leaf_net283;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net262;
 wire clknet_1_0__leaf_net262;
 wire clknet_1_1__leaf_net262;
 wire clknet_0_net251;
 wire clknet_1_0__leaf_net251;
 wire clknet_1_1__leaf_net251;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net701;
 wire clknet_1_0__leaf_net701;
 wire clknet_1_1__leaf_net701;
 wire clknet_0_net258;
 wire clknet_1_0__leaf_net258;
 wire clknet_1_1__leaf_net258;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net244;
 wire clknet_1_0__leaf_net244;
 wire clknet_1_1__leaf_net244;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;

 sky130_fd_sc_hd__a41o_2 c100 (.A1(net33),
    .A2(net21),
    .A3(net35),
    .A4(net36),
    .B1(net956),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c101 (.A0(net938),
    .A1(net28),
    .A2(net35),
    .A3(net847),
    .S0(net36),
    .S1(net33),
    .X(net38));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net32),
    .A2(net36),
    .B1_N(net987),
    .X(net39));
 sky130_fd_sc_hd__mux4_1 c103 (.A0(net38),
    .A1(net5),
    .A2(net37),
    .A3(net33),
    .S0(net28),
    .S1(net35),
    .X(net40));
 sky130_fd_sc_hd__xnor2_2 c104 (.A(net34),
    .B(net824),
    .Y(net41));
 sky130_fd_sc_hd__a41o_2 c105 (.A1(net30),
    .A2(net37),
    .A3(net41),
    .A4(net31),
    .B1(net33),
    .X(net42));
 sky130_fd_sc_hd__xnor2_1 c106 (.A(net35),
    .B(net36),
    .Y(net43));
 sky130_fd_sc_hd__a21bo_1 c107 (.A1(net43),
    .A2(net31),
    .B1_N(net41),
    .X(net44));
 sky130_fd_sc_hd__a41o_1 c108 (.A1(net39),
    .A2(net43),
    .A3(net44),
    .A4(net31),
    .B1(net30),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net44),
    .A1(net33),
    .A2(net9),
    .A3(net983),
    .S0(net42),
    .S1(net34),
    .X(net46));
 sky130_fd_sc_hd__xnor2_4 c110 (.A(net856),
    .B(net876),
    .Y(net47));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net847),
    .B(net31),
    .Y(net48));
 sky130_fd_sc_hd__a21bo_2 c112 (.A1(net873),
    .A2(net944),
    .B1_N(net847),
    .X(net49));
 sky130_fd_sc_hd__xnor2_1 c113 (.A(net49),
    .B(net944),
    .Y(net50));
 sky130_fd_sc_hd__xnor2_1 c114 (.A(net47),
    .B(net49),
    .Y(net51));
 sky130_fd_sc_hd__clkbuf_1 c115 (.A(net679),
    .X(net52));
 sky130_fd_sc_hd__xnor2_2 c116 (.A(net47),
    .B(net49),
    .Y(net914));
 sky130_fd_sc_hd__xnor2_1 c117 (.A(net31),
    .B(net36),
    .Y(net53));
 sky130_fd_sc_hd__clkbuf_1 c118 (.A(net679),
    .X(net54));
 sky130_fd_sc_hd__a21bo_1 c119 (.A1(net48),
    .A2(net52),
    .B1_N(net36),
    .X(net55));
 sky130_fd_sc_hd__a21bo_1 c120 (.A1(net36),
    .A2(net47),
    .B1_N(net944),
    .X(net56));
 sky130_fd_sc_hd__xnor2_2 c121 (.A(net854),
    .B(net944),
    .Y(net921));
 sky130_fd_sc_hd__mux4_1 c122 (.A0(net55),
    .A1(net26),
    .A2(net31),
    .A3(net56),
    .S0(net48),
    .S1(net921),
    .X(net57));
 sky130_fd_sc_hd__buf_1 c123 (.A(net728),
    .X(net926));
 sky130_fd_sc_hd__a31o_1 c124 (.A1(net53),
    .A2(net921),
    .A3(net926),
    .B1(net47),
    .X(net58));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net57),
    .A1(net49),
    .A2(net46),
    .A3(net36),
    .S0(net31),
    .S1(net53),
    .X(net59));
 sky130_fd_sc_hd__a21bo_1 c126 (.A1(net26),
    .A2(net56),
    .B1_N(net921),
    .X(net60));
 sky130_fd_sc_hd__buf_1 c127 (.A(net678),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 c128 (.A(net728),
    .X(net916));
 sky130_fd_sc_hd__a21bo_2 c129 (.A1(net52),
    .A2(net916),
    .B1_N(net56),
    .X(net928));
 sky130_fd_sc_hd__sdfrbp_1 c130 (.CLK(clknet_4_10_0_clk),
    .D(net869),
    .RESET_B(net928),
    .SCD(net37),
    .SCE(net60),
    .Q(net881),
    .Q_N(net62));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net60),
    .A1(net928),
    .A2(net61),
    .A3(net62),
    .S0(net37),
    .S1(net55),
    .X(net63));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net618),
    .B(net874),
    .Y(net64));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net825),
    .B(net820),
    .Y(net65));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net819),
    .B(net826),
    .Y(net66));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net671),
    .B(net820),
    .Y(net67));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net66),
    .B(net822),
    .Y(net68));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net65),
    .B(net838),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_4 c138 (.A(net68),
    .B(net874),
    .Y(net887));
 sky130_fd_sc_hd__xnor2_2 c139 (.A(net887),
    .B(net968),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_4 c140 (.A(net69),
    .B(net838),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_4 c141 (.A(net66),
    .B(net961),
    .Y(net72));
 sky130_fd_sc_hd__a21bo_2 c142 (.A1(net874),
    .A2(net72),
    .B1_N(net860),
    .X(net73));
 sky130_fd_sc_hd__xnor2_2 c143 (.A(net817),
    .B(net849),
    .Y(net74));
 sky130_fd_sc_hd__xnor2_4 c144 (.A(net72),
    .B(net819),
    .Y(net75));
 sky130_fd_sc_hd__xnor2_4 c145 (.A(net64),
    .B(net72),
    .Y(net76));
 sky130_fd_sc_hd__a21bo_1 c146 (.A1(net824),
    .A2(net825),
    .B1_N(net820),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net820),
    .A1(net75),
    .A2(net77),
    .A3(net66),
    .S0(net71),
    .S1(net67),
    .X(net78));
 sky130_fd_sc_hd__a31o_4 c148 (.A1(net65),
    .A2(net76),
    .A3(net78),
    .B1(net73),
    .X(net79));
 sky130_fd_sc_hd__a41o_4 c149 (.A1(net826),
    .A2(net76),
    .A3(net77),
    .A4(net959),
    .B1(net65),
    .X(net80));
 sky130_fd_sc_hd__a21bo_2 c150 (.A1(net77),
    .A2(net73),
    .B1_N(net79),
    .X(net81));
 sky130_fd_sc_hd__a31o_4 c151 (.A1(net73),
    .A2(net71),
    .A3(net81),
    .B1(net79),
    .X(net82));
 sky130_fd_sc_hd__xnor2_4 c152 (.A(net71),
    .B(net81),
    .Y(net83));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net838),
    .A1(net80),
    .A2(net83),
    .A3(net849),
    .S0(net81),
    .S1(net82),
    .X(net84));
 sky130_fd_sc_hd__xnor2_1 c154 (.A(net83),
    .B(net875),
    .Y(net85));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net967),
    .B(net83),
    .Y(net878));
 sky130_fd_sc_hd__xnor2_2 c156 (.A(net839),
    .B(net821),
    .Y(net86));
 sky130_fd_sc_hd__a31o_1 c157 (.A1(net85),
    .A2(net67),
    .A3(net959),
    .B1(net84),
    .X(net87));
 sky130_fd_sc_hd__a21bo_4 c158 (.A1(net841),
    .A2(net849),
    .B1_N(net950),
    .X(net88));
 sky130_fd_sc_hd__a21bo_2 c159 (.A1(net850),
    .A2(net949),
    .B1_N(net831),
    .X(net89));
 sky130_fd_sc_hd__a31o_1 c160 (.A1(net846),
    .A2(net89),
    .A3(net853),
    .B1(net949),
    .X(net90));
 sky130_fd_sc_hd__a21bo_4 c161 (.A1(net848),
    .A2(net949),
    .B1_N(net831),
    .X(net91));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net949),
    .B(net953),
    .Y(net92));
 sky130_fd_sc_hd__a21bo_1 c163 (.A1(net843),
    .A2(net92),
    .B1_N(net949),
    .X(net93));
 sky130_fd_sc_hd__a21bo_4 c164 (.A1(net853),
    .A2(net93),
    .B1_N(net91),
    .X(net94));
 sky130_fd_sc_hd__a21bo_4 c165 (.A1(net92),
    .A2(net83),
    .B1_N(net88),
    .X(net95));
 sky130_fd_sc_hd__a21bo_1 c166 (.A1(net90),
    .A2(net92),
    .B1_N(net94),
    .X(net96));
 sky130_fd_sc_hd__a21bo_1 c167 (.A1(net837),
    .A2(net851),
    .B1_N(net949),
    .X(net97));
 sky130_fd_sc_hd__a21bo_1 c168 (.A1(net849),
    .A2(net848),
    .B1_N(net949),
    .X(net98));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net98),
    .A1(net97),
    .A2(net86),
    .A3(net92),
    .S0(net959),
    .S1(net836),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 c170 (.A0(net96),
    .A1(net850),
    .A2(net97),
    .A3(net92),
    .S0(net99),
    .S1(net85),
    .X(net100));
 sky130_fd_sc_hd__buf_1 c171 (.A(net692),
    .X(net101));
 sky130_fd_sc_hd__a21bo_1 c172 (.A1(net97),
    .A2(net949),
    .B1_N(net99),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 c173 (.A(net692),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c174 (.A0(net103),
    .A1(net85),
    .A2(net100),
    .A3(net102),
    .S0(net89),
    .S1(net88),
    .X(net104));
 sky130_fd_sc_hd__mux4_2 c175 (.A0(net89),
    .A1(net96),
    .A2(net103),
    .A3(net101),
    .S0(net959),
    .S1(net845),
    .X(net105));
 sky130_fd_sc_hd__a21bo_1 c176 (.A1(net67),
    .A2(net94),
    .B1_N(net76),
    .X(net106));
 sky130_fd_sc_hd__xnor2_2 c177 (.A(net99),
    .B(net865),
    .Y(net107));
 sky130_fd_sc_hd__xnor2_1 c178 (.A(net107),
    .B(net828),
    .Y(net108));
 sky130_fd_sc_hd__xnor2_2 c179 (.A(net844),
    .B(net862),
    .Y(net109));
 sky130_fd_sc_hd__a21bo_1 c180 (.A1(net840),
    .A2(net855),
    .B1_N(net94),
    .X(net110));
 sky130_fd_sc_hd__a21bo_1 c181 (.A1(net110),
    .A2(net109),
    .B1_N(net950),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 c182 (.A(net668),
    .X(net112));
 sky130_fd_sc_hd__a31o_1 c183 (.A1(net90),
    .A2(net67),
    .A3(net110),
    .B1(net953),
    .X(net113));
 sky130_fd_sc_hd__xnor2_2 c184 (.A(net832),
    .B(net863),
    .Y(net114));
 sky130_fd_sc_hd__a21bo_2 c185 (.A1(net3),
    .A2(net94),
    .B1_N(net854),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 c186 (.A(net668),
    .X(net116));
 sky130_fd_sc_hd__a21bo_1 c187 (.A1(net114),
    .A2(net953),
    .B1_N(net943),
    .X(net117));
 sky130_fd_sc_hd__a41o_1 c188 (.A1(net113),
    .A2(net109),
    .A3(net943),
    .A4(net107),
    .B1(net830),
    .X(net118));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net868),
    .A1(net107),
    .A2(net861),
    .A3(net84),
    .S0(net943),
    .S1(net717),
    .X(net119));
 sky130_fd_sc_hd__a31o_1 c190 (.A1(net119),
    .A2(net107),
    .A3(net94),
    .X(net120));
 sky130_fd_sc_hd__sdfrbp_1 c191 (.CLK(clknet_4_2_0_clk),
    .D(net108),
    .RESET_B(net73),
    .SCD(net851),
    .SCE(net111),
    .Q(net122),
    .Q_N(net121));
 sky130_fd_sc_hd__a41o_4 c192 (.A1(net943),
    .A2(net114),
    .A3(net90),
    .A4(net950),
    .B1(net717),
    .X(net123));
 sky130_fd_sc_hd__sdfrtn_1 c193 (.CLK_N(clknet_4_2_0_clk),
    .D(net116),
    .RESET_B(net113),
    .SCD(net117),
    .SCE(net717),
    .Q(net124));
 sky130_fd_sc_hd__a31o_2 c194 (.A1(net109),
    .A2(net122),
    .A3(net968),
    .B1(net717),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net111),
    .A1(net124),
    .A2(net125),
    .A3(net121),
    .S0(net123),
    .S1(net717),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 c196 (.A(net668),
    .X(net127));
 sky130_fd_sc_hd__a41o_4 c197 (.A1(net127),
    .A2(net122),
    .A3(net114),
    .A4(net124),
    .B1(net717),
    .X(net128));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net16),
    .A2(net23),
    .B1_N(net995),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net972),
    .A1(net845),
    .A2(net88),
    .A3(net975),
    .S0(net75),
    .S1(net980),
    .X(net130));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net19),
    .A2(net20),
    .B1_N(net970),
    .X(net131));
 sky130_fd_sc_hd__xnor2_4 c201 (.A(net129),
    .B(net944),
    .Y(net132));
 sky130_fd_sc_hd__a21bo_2 c202 (.A1(net17),
    .A2(net125),
    .B1_N(net692),
    .X(net133));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net124),
    .A2(net971),
    .B1_N(net112),
    .X(net134));
 sky130_fd_sc_hd__a21bo_2 c204 (.A1(net134),
    .A2(net132),
    .B1_N(net951),
    .X(net135));
 sky130_fd_sc_hd__a41o_1 c205 (.A1(net130),
    .A2(net135),
    .A3(net84),
    .A4(net132),
    .B1(net17),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 c206 (.A(net1017),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 c207 (.A(net708),
    .X(net138));
 sky130_fd_sc_hd__sdfbbn_2 c208 (.CLK_N(clknet_4_8_0_clk),
    .D(net135),
    .RESET_B(net863),
    .SCD(net132),
    .SCE(net11),
    .SET_B(net128),
    .Q(net140),
    .Q_N(net139));
 sky130_fd_sc_hd__a31o_2 c209 (.A1(net91),
    .A2(net132),
    .A3(net955),
    .B1(net692),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net141),
    .A1(net128),
    .A2(net976),
    .A3(net944),
    .S0(net950),
    .S1(net7),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 c211 (.A(net668),
    .X(net913));
 sky130_fd_sc_hd__sdfrtp_4 c212 (.CLK(clknet_4_8_0_clk),
    .D(net138),
    .RESET_B(net960),
    .SCD(net141),
    .SCE(net740),
    .Q(net929));
 sky130_fd_sc_hd__mux4_1 c213 (.A0(net7),
    .A1(net135),
    .A2(net835),
    .A3(net929),
    .S0(net997),
    .S1(net740),
    .X(net143));
 sky130_fd_sc_hd__a41o_1 c214 (.A1(net137),
    .A2(net960),
    .A3(net132),
    .A4(net692),
    .B1(net964),
    .X(net144));
 sky130_fd_sc_hd__a31o_1 c215 (.A1(net141),
    .A2(net960),
    .A3(net943),
    .B1(net715),
    .X(net145));
 sky130_fd_sc_hd__sdfbbn_1 c216 (.CLK_N(clknet_4_8_0_clk),
    .D(net845),
    .RESET_B(net140),
    .SCD(net117),
    .SCE(net929),
    .SET_B(net141),
    .Q(net147),
    .Q_N(net146));
 sky130_fd_sc_hd__a31o_1 c217 (.A1(net147),
    .A2(net95),
    .A3(net960),
    .B1(net715),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net117),
    .A1(net148),
    .A2(net959),
    .A3(net123),
    .S0(net740),
    .S1(net964),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net117),
    .A1(net146),
    .A2(net148),
    .A3(net135),
    .S0(net929),
    .S1(net714),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 c220 (.A(net708),
    .X(net151));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(net128),
    .B(net115),
    .Y(net152));
 sky130_fd_sc_hd__xnor2_4 c222 (.A(net32),
    .B(net824),
    .Y(net153));
 sky130_fd_sc_hd__xnor2_4 c223 (.A(net140),
    .B(net128),
    .Y(net880));
 sky130_fd_sc_hd__a21bo_1 c224 (.A1(net73),
    .A2(net978),
    .B1_N(net964),
    .X(net154));
 sky130_fd_sc_hd__xnor2_2 c225 (.A(net11),
    .B(net42),
    .Y(net155));
 sky130_fd_sc_hd__a41o_1 c226 (.A1(net141),
    .A2(net128),
    .A3(net42),
    .A4(net148),
    .B1(net938),
    .X(net156));
 sky130_fd_sc_hd__xnor2_4 c227 (.A(net153),
    .B(net95),
    .Y(net893));
 sky130_fd_sc_hd__mux4_1 c228 (.A0(net155),
    .A1(net5),
    .A2(net154),
    .A3(net135),
    .S0(net42),
    .S1(net964),
    .X(net157));
 sky130_fd_sc_hd__a21bo_1 c229 (.A1(net132),
    .A2(net865),
    .B1_N(clknet_1_0__leaf_net743),
    .X(net158));
 sky130_fd_sc_hd__xnor2_2 c230 (.A(net153),
    .B(net929),
    .Y(net923));
 sky130_fd_sc_hd__buf_1 c231 (.A(net670),
    .X(net159));
 sky130_fd_sc_hd__buf_1 c232 (.A(net670),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 c233 (.A0(net1),
    .A1(net159),
    .A2(net155),
    .A3(net880),
    .S0(net132),
    .S1(net33),
    .X(net161));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net42),
    .A2(net893),
    .B1_N(clknet_1_0__leaf_net743),
    .X(net162));
 sky130_fd_sc_hd__buf_1 c235 (.A(net708),
    .X(net918));
 sky130_fd_sc_hd__mux4_1 c236 (.A0(clknet_1_1__leaf_net158),
    .A1(clknet_1_0__leaf_net162),
    .A2(net32),
    .A3(net938),
    .S0(net960),
    .S1(net42),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c237 (.A0(net5),
    .A1(net11),
    .A2(net45),
    .A3(net161),
    .S0(net938),
    .S1(net153),
    .X(net164));
 sky130_fd_sc_hd__xnor2_1 c238 (.A(clknet_1_1__leaf_net162),
    .B(net745),
    .Y(net165));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net923),
    .A1(net91),
    .A2(net144),
    .A3(net141),
    .S0(net155),
    .S1(net744),
    .X(net166));
 sky130_fd_sc_hd__sdfbbp_1 c240 (.CLK(clknet_4_10_0_clk),
    .D(net161),
    .RESET_B(clknet_1_0__leaf_net165),
    .SCD(net992),
    .SCE(clknet_1_1__leaf_net743),
    .SET_B(net744),
    .Q(net168),
    .Q_N(net167));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_1__leaf_net165),
    .A1(net938),
    .A2(net160),
    .A3(net168),
    .S0(net880),
    .S1(clknet_1_1__leaf_net743),
    .X(net169));
 sky130_fd_sc_hd__sdfrtp_1 c242 (.CLK(clknet_4_10_0_clk),
    .D(net943),
    .RESET_B(net914),
    .SCD(net37),
    .SCE(net964),
    .Q(net931));
 sky130_fd_sc_hd__a21bo_1 c243 (.A1(net37),
    .A2(net840),
    .B1_N(net944),
    .X(net925));
 sky130_fd_sc_hd__a21bo_1 c244 (.A1(net929),
    .A2(net41),
    .B1_N(net736),
    .X(net170));
 sky130_fd_sc_hd__a41o_1 c245 (.A1(net56),
    .A2(net916),
    .A3(net840),
    .A4(net943),
    .B1(net737),
    .X(net171));
 sky130_fd_sc_hd__a21bo_1 c246 (.A1(net840),
    .A2(net943),
    .B1_N(net37),
    .X(net896));
 sky130_fd_sc_hd__buf_1 c247 (.A(net728),
    .X(net172));
 sky130_fd_sc_hd__a21bo_1 c248 (.A1(net172),
    .A2(net893),
    .B1_N(net37),
    .X(net173));
 sky130_fd_sc_hd__xnor2_1 c249 (.A(net45),
    .B(net172),
    .Y(net174));
 sky130_fd_sc_hd__a21bo_1 c250 (.A1(net943),
    .A2(net840),
    .B1_N(net855),
    .X(net917));
 sky130_fd_sc_hd__buf_1 c251 (.A(net728),
    .X(net175));
 sky130_fd_sc_hd__a21bo_1 c252 (.A1(net855),
    .A2(net175),
    .B1_N(net931),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net174),
    .A1(net172),
    .A2(net893),
    .A3(net960),
    .S0(net175),
    .S1(net171),
    .X(net177));
 sky130_fd_sc_hd__a31o_1 c254 (.A1(net58),
    .A2(net736),
    .A3(net738),
    .B1(net748),
    .X(net178));
 sky130_fd_sc_hd__a41o_1 c255 (.A1(net923),
    .A2(net175),
    .A3(net62),
    .A4(net735),
    .B1(net748),
    .X(net904));
 sky130_fd_sc_hd__a21bo_1 c256 (.A1(net925),
    .A2(net745),
    .B1_N(net746),
    .X(net934));
 sky130_fd_sc_hd__a21bo_1 c257 (.A1(net41),
    .A2(net115),
    .B1_N(net670),
    .X(net915));
 sky130_fd_sc_hd__buf_1 c258 (.A(net678),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net175),
    .A1(net37),
    .A2(net172),
    .A3(net931),
    .S0(net934),
    .S1(net738),
    .X(net180));
 sky130_fd_sc_hd__mux4_2 c260 (.A0(net173),
    .A1(net172),
    .A2(net175),
    .A3(net881),
    .S0(net179),
    .S1(net748),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c261 (.A0(net176),
    .A1(net179),
    .A2(net895),
    .A3(net893),
    .S0(net735),
    .S1(net748),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net895),
    .A1(net914),
    .A2(net931),
    .A3(net670),
    .S0(clknet_1_1__leaf_net919),
    .S1(net748),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net61),
    .A1(net931),
    .A2(net895),
    .A3(clknet_1_0__leaf_net891),
    .S0(clknet_1_0__leaf_net919),
    .S1(net903),
    .X(net183));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net828),
    .B(net78),
    .Y(net184));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net80),
    .B(net967),
    .Y(net185));
 sky130_fd_sc_hd__xnor2_2 c266 (.A(net818),
    .B(net78),
    .Y(net186));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net79),
    .B(net80),
    .Y(net187));
 sky130_fd_sc_hd__xnor2_4 c268 (.A(net68),
    .B(net184),
    .Y(net188));
 sky130_fd_sc_hd__xnor2_1 c269 (.A(net829),
    .B(net188),
    .Y(net189));
 sky130_fd_sc_hd__xnor2_1 c270 (.A(net78),
    .B(net186),
    .Y(net190));
 sky130_fd_sc_hd__xnor2_1 c271 (.A(net188),
    .B(net187),
    .Y(net191));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net823),
    .B(net79),
    .Y(net192));
 sky130_fd_sc_hd__a21bo_1 c273 (.A1(net187),
    .A2(net184),
    .B1_N(net186),
    .X(net193));
 sky130_fd_sc_hd__a21bo_1 c274 (.A1(net191),
    .A2(net193),
    .B1_N(net75),
    .X(net194));
 sky130_fd_sc_hd__a21bo_2 c275 (.A1(net189),
    .A2(net959),
    .B1_N(net186),
    .X(net195));
 sky130_fd_sc_hd__mux4_1 c276 (.A0(net185),
    .A1(net78),
    .A2(net186),
    .A3(net68),
    .S0(net195),
    .S1(net959),
    .X(net196));
 sky130_fd_sc_hd__a21bo_2 c277 (.A1(net79),
    .A2(net78),
    .B1_N(net196),
    .X(net197));
 sky130_fd_sc_hd__a21bo_1 c278 (.A1(net191),
    .A2(net189),
    .B1_N(net195),
    .X(net198));
 sky130_fd_sc_hd__a31o_2 c279 (.A1(net184),
    .A2(net197),
    .A3(net192),
    .B1(net188),
    .X(net199));
 sky130_fd_sc_hd__a21bo_1 c280 (.A1(net196),
    .A2(net198),
    .B1_N(net199),
    .X(net930));
 sky130_fd_sc_hd__a21bo_2 c281 (.A1(net198),
    .A2(net947),
    .B1_N(net189),
    .X(net200));
 sky130_fd_sc_hd__a21bo_1 c282 (.A1(net186),
    .A2(net199),
    .B1_N(net194),
    .X(net201));
 sky130_fd_sc_hd__a31o_2 c283 (.A1(net194),
    .A2(net199),
    .A3(net196),
    .B1(net947),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net946),
    .A1(net200),
    .A2(net190),
    .A3(net194),
    .S0(net195),
    .S1(net198),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net203),
    .A1(net191),
    .A2(net946),
    .A3(net194),
    .S0(net947),
    .S1(net202),
    .X(net204));
 sky130_fd_sc_hd__a21bo_1 c286 (.A1(net89),
    .A2(net875),
    .B1_N(net190),
    .X(net205));
 sky130_fd_sc_hd__a21bo_1 c287 (.A1(net101),
    .A2(net195),
    .B1_N(net949),
    .X(net206));
 sky130_fd_sc_hd__a21bo_4 c288 (.A1(net205),
    .A2(net202),
    .B1_N(net851),
    .X(net207));
 sky130_fd_sc_hd__a21bo_4 c289 (.A1(net851),
    .A2(net953),
    .B1_N(net842),
    .X(net208));
 sky130_fd_sc_hd__a21bo_1 c290 (.A1(net875),
    .A2(net101),
    .B1_N(net208),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c291 (.A0(net207),
    .A1(net76),
    .A2(net195),
    .A3(net860),
    .S0(net937),
    .S1(net91),
    .X(net210));
 sky130_fd_sc_hd__a21bo_1 c292 (.A1(net98),
    .A2(net94),
    .B1_N(net92),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net209),
    .A1(net192),
    .A2(net207),
    .A3(net185),
    .S0(net208),
    .S1(net202),
    .X(net212));
 sky130_fd_sc_hd__a21bo_1 c294 (.A1(net205),
    .A2(net95),
    .B1_N(net93),
    .X(net213));
 sky130_fd_sc_hd__a21bo_1 c295 (.A1(net101),
    .A2(net88),
    .B1_N(net750),
    .X(net214));
 sky130_fd_sc_hd__a31o_1 c296 (.A1(net190),
    .A2(net211),
    .A3(net199),
    .B1(net950),
    .X(net215));
 sky130_fd_sc_hd__a21bo_2 c297 (.A1(net209),
    .A2(net669),
    .B1_N(net750),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 c298 (.A(net669),
    .X(net217));
 sky130_fd_sc_hd__a41o_1 c299 (.A1(net211),
    .A2(net946),
    .A3(net216),
    .A4(net215),
    .B1(net950),
    .X(net218));
 sky130_fd_sc_hd__mux4_2 c300 (.A0(net214),
    .A1(net216),
    .A2(net209),
    .A3(net91),
    .S0(net946),
    .S1(net206),
    .X(net219));
 sky130_fd_sc_hd__a21bo_1 c301 (.A1(net89),
    .A2(net217),
    .B1_N(net750),
    .X(net220));
 sky130_fd_sc_hd__mux4_2 c302 (.A0(net93),
    .A1(net206),
    .A2(net209),
    .A3(net91),
    .S0(net711),
    .S1(net749),
    .X(net221));
 sky130_fd_sc_hd__mux4_2 c303 (.A0(net217),
    .A1(net831),
    .A2(net213),
    .A3(net221),
    .S0(net219),
    .S1(net711),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 c304 (.A(net669),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net223),
    .A1(net220),
    .A2(net222),
    .A3(net213),
    .S0(net202),
    .X(net224));
 sky130_fd_sc_hd__a41o_2 c306 (.A1(net206),
    .A2(net75),
    .A3(net208),
    .A4(net221),
    .B1(net711),
    .X(net892));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net219),
    .A1(net89),
    .A2(net211),
    .A3(net222),
    .S0(net207),
    .S1(net711),
    .X(net225));
 sky130_fd_sc_hd__xnor2_2 c308 (.A(net94),
    .B(net739),
    .Y(net226));
 sky130_fd_sc_hd__xnor2_2 c309 (.A(net830),
    .B(net82),
    .Y(net227));
 sky130_fd_sc_hd__a21bo_1 c310 (.A1(net102),
    .A2(net125),
    .B1_N(net750),
    .X(net228));
 sky130_fd_sc_hd__xnor2_2 c311 (.A(net858),
    .B(net213),
    .Y(net229));
 sky130_fd_sc_hd__xnor2_1 c312 (.A(net202),
    .B(net711),
    .Y(net230));
 sky130_fd_sc_hd__xnor2_4 c313 (.A(net216),
    .B(net952),
    .Y(net231));
 sky130_fd_sc_hd__a41o_1 c314 (.A1(net213),
    .A2(net112),
    .A3(net947),
    .A4(net937),
    .B1(net123),
    .X(net232));
 sky130_fd_sc_hd__sdfrtp_1 c315 (.CLK(clknet_4_2_0_clk),
    .D(net842),
    .RESET_B(net950),
    .SCD(net119),
    .SCE(net208),
    .Q(net233));
 sky130_fd_sc_hd__a41o_1 c316 (.A1(net0),
    .A2(net102),
    .A3(net952),
    .A4(net125),
    .B1(net119),
    .X(net234));
 sky130_fd_sc_hd__a21bo_2 c317 (.A1(net221),
    .A2(net947),
    .B1_N(net687),
    .X(net235));
 sky130_fd_sc_hd__mux4_2 c318 (.A0(net202),
    .A1(net832),
    .A2(net82),
    .A3(net231),
    .S0(net851),
    .S1(net233),
    .X(net236));
 sky130_fd_sc_hd__a21bo_1 c319 (.A1(net233),
    .A2(net216),
    .B1_N(net687),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net195),
    .A1(net123),
    .A2(net124),
    .A3(net125),
    .S0(net952),
    .S1(net854),
    .X(net238));
 sky130_fd_sc_hd__xnor2_2 c321 (.A(net226),
    .B(net739),
    .Y(net239));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net237),
    .A2(net942),
    .B1_N(net235),
    .X(net240));
 sky130_fd_sc_hd__a21bo_1 c323 (.A1(net199),
    .A2(net228),
    .B1_N(net231),
    .X(net241));
 sky130_fd_sc_hd__mux4_2 c324 (.A0(net211),
    .A1(net235),
    .A2(net226),
    .A3(net942),
    .S0(net228),
    .S1(net739),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net236),
    .A1(net241),
    .A2(net240),
    .A3(net231),
    .S0(net739),
    .S1(net752),
    .X(net243));
 sky130_fd_sc_hd__a41o_1 c326 (.A1(net219),
    .A2(net124),
    .A3(net102),
    .A4(clknet_1_0__leaf_net701),
    .B1(net753),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(clknet_1_0__leaf_net244),
    .A1(net237),
    .A2(net242),
    .A3(net952),
    .S0(clknet_1_0__leaf_net701),
    .S1(net752),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net240),
    .A1(net236),
    .A2(clknet_1_1__leaf_net244),
    .A3(net952),
    .S0(net752),
    .S1(net754),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net235),
    .A1(net240),
    .A2(net937),
    .A3(net753),
    .S0(net755),
    .S1(net756),
    .X(net247));
 sky130_fd_sc_hd__xnor2_2 c330 (.A(net980),
    .B(net124),
    .Y(net248));
 sky130_fd_sc_hd__a21bo_1 c331 (.A1(net929),
    .A2(net964),
    .B1_N(clknet_1_1__leaf_net742),
    .X(net249));
 sky130_fd_sc_hd__a41o_1 c332 (.A1(net208),
    .A2(net123),
    .A3(net197),
    .A4(net851),
    .B1(net124),
    .X(net250));
 sky130_fd_sc_hd__a21bo_1 c333 (.A1(net249),
    .A2(net946),
    .B1_N(net929),
    .X(net251));
 sky130_fd_sc_hd__a21bo_1 c334 (.A1(net124),
    .A2(net955),
    .B1_N(net687),
    .X(net908));
 sky130_fd_sc_hd__buf_1 c335 (.A(net726),
    .X(net252));
 sky130_fd_sc_hd__a21bo_2 c336 (.A1(net112),
    .A2(net139),
    .B1_N(net753),
    .X(net253));
 sky130_fd_sc_hd__a21bo_1 c337 (.A1(net681),
    .A2(net687),
    .B1_N(clknet_1_1__leaf_net701),
    .X(net902));
 sky130_fd_sc_hd__a41o_1 c338 (.A1(net252),
    .A2(net867),
    .A3(net84),
    .A4(net942),
    .B1(net112),
    .X(net254));
 sky130_fd_sc_hd__a31o_1 c339 (.A1(net233),
    .A2(net948),
    .A3(net988),
    .B1(clknet_1_0__leaf_net742),
    .X(net255));
 sky130_fd_sc_hd__a21bo_1 c340 (.A1(net975),
    .A2(net248),
    .B1_N(clknet_1_0__leaf_net742),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net207),
    .A1(net969),
    .A2(net230),
    .A3(net835),
    .S0(net937),
    .S1(net1009),
    .X(net257));
 sky130_fd_sc_hd__a41o_1 c342 (.A1(net140),
    .A2(net851),
    .A3(net253),
    .A4(clknet_1_1__leaf_net701),
    .B1(net753),
    .X(net258));
 sky130_fd_sc_hd__sdfbbn_2 c343 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net258),
    .RESET_B(net254),
    .SCD(clknet_1_0__leaf_net251),
    .SCE(net253),
    .SET_B(net981),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__a41o_1 c344 (.A1(net84),
    .A2(net223),
    .A3(clknet_1_1__leaf_net902),
    .A4(net823),
    .B1(clknet_1_0__leaf_net251),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c345 (.A0(net147),
    .A1(net253),
    .A2(net124),
    .A3(clknet_1_0__leaf_net255),
    .S0(clknet_1_0__leaf_net251),
    .S1(net680),
    .X(net262));
 sky130_fd_sc_hd__buf_2 c346 (.A(net726),
    .X(net263));
 sky130_fd_sc_hd__a41o_1 c347 (.A1(clknet_1_1__leaf_net258),
    .A2(net263),
    .A3(clknet_1_0__leaf_net251),
    .A4(clknet_1_1__leaf_net261),
    .B1(net123),
    .X(net264));
 sky130_fd_sc_hd__a41o_2 c348 (.A1(net988),
    .A2(net263),
    .A3(net253),
    .A4(net680),
    .B1(net898),
    .X(net905));
 sky130_fd_sc_hd__a41o_1 c349 (.A1(clknet_1_0__leaf_net261),
    .A2(net905),
    .A3(net259),
    .A4(clknet_1_0__leaf_net251),
    .B1(net835),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 c350 (.A(net727),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net266),
    .A1(clknet_1_0__leaf_net261),
    .A2(net146),
    .A3(net254),
    .S0(net208),
    .S1(net898),
    .X(net267));
 sky130_fd_sc_hd__buf_1 c352 (.A(net675),
    .X(net268));
 sky130_fd_sc_hd__buf_2 c353 (.A(net675),
    .X(net269));
 sky130_fd_sc_hd__a21bo_2 c354 (.A1(net269),
    .A2(net978),
    .B1_N(net757),
    .X(net270));
 sky130_fd_sc_hd__xnor2_1 c355 (.A(net154),
    .B(net269),
    .Y(net271));
 sky130_fd_sc_hd__xnor2_1 c356 (.A(net132),
    .B(net263),
    .Y(net272));
 sky130_fd_sc_hd__xnor2_1 c357 (.A(net160),
    .B(net749),
    .Y(net273));
 sky130_fd_sc_hd__buf_1 c358 (.A(net727),
    .X(net274));
 sky130_fd_sc_hd__xnor2_1 c359 (.A(net95),
    .B(net932),
    .Y(net275));
 sky130_fd_sc_hd__a21bo_1 c360 (.A1(net271),
    .A2(net269),
    .B1_N(net867),
    .X(net276));
 sky130_fd_sc_hd__xnor2_1 c361 (.A(net274),
    .B(net270),
    .Y(net277));
 sky130_fd_sc_hd__a21bo_2 c362 (.A1(net275),
    .A2(net273),
    .B1_N(net747),
    .X(net897));
 sky130_fd_sc_hd__xnor2_1 c363 (.A(net273),
    .B(net277),
    .Y(net278));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net970),
    .A1(net905),
    .A2(net897),
    .A3(net274),
    .S0(net269),
    .S1(net254),
    .X(net279));
 sky130_fd_sc_hd__a21bo_1 c365 (.A1(net33),
    .A2(clknet_1_1__leaf_net251),
    .B1_N(net758),
    .X(net280));
 sky130_fd_sc_hd__xnor2_1 c366 (.A(net252),
    .B(net269),
    .Y(net281));
 sky130_fd_sc_hd__a21bo_1 c367 (.A1(net33),
    .A2(net268),
    .B1_N(net758),
    .X(net922));
 sky130_fd_sc_hd__xnor2_1 c368 (.A(net268),
    .B(net948),
    .Y(net282));
 sky130_fd_sc_hd__a21bo_1 c369 (.A1(net282),
    .A2(clknet_1_0__leaf_net256),
    .B1_N(net758),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net148),
    .A1(net128),
    .A2(net281),
    .A3(net897),
    .S0(net275),
    .S1(net758),
    .X(net284));
 sky130_fd_sc_hd__a21bo_2 c371 (.A1(net277),
    .A2(net269),
    .B1_N(net988),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net284),
    .A1(net893),
    .A2(net897),
    .A3(net285),
    .S0(net167),
    .S1(net758),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net281),
    .A1(net282),
    .A2(net263),
    .A3(net984),
    .S0(net675),
    .S1(net758),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net280),
    .A1(net75),
    .A2(net918),
    .A3(net914),
    .S0(net928),
    .S1(net916),
    .X(net288));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net287),
    .A1(net892),
    .A2(net918),
    .A3(net681),
    .S0(net964),
    .S1(clknet_1_0__leaf_net906),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net91),
    .A1(net61),
    .A2(net926),
    .A3(net892),
    .S0(net925),
    .S1(net903),
    .X(net884));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(clknet_1_1__leaf_net255),
    .A1(net287),
    .A3(clknet_1_0__leaf_net891),
    .S0(net903),
    .S1(clknet_1_0__leaf_net906),
    .X(net290));
 sky130_fd_sc_hd__xnor2_4 c396 (.A(net84),
    .B(net188),
    .Y(net291));
 sky130_fd_sc_hd__a21bo_2 c397 (.A1(net188),
    .A2(net291),
    .B1_N(net84),
    .X(net292));
 sky130_fd_sc_hd__a21bo_1 c398 (.A1(net291),
    .A2(net192),
    .B1_N(net947),
    .X(net293));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net822),
    .B(net185),
    .Y(net294));
 sky130_fd_sc_hd__a21bo_1 c400 (.A1(net193),
    .A2(net84),
    .B1_N(net293),
    .X(net295));
 sky130_fd_sc_hd__buf_2 c401 (.A(net664),
    .X(net879));
 sky130_fd_sc_hd__a21bo_1 c402 (.A1(net293),
    .A2(net821),
    .B1_N(net70),
    .X(net296));
 sky130_fd_sc_hd__a21bo_1 c403 (.A1(net671),
    .A2(net871),
    .B1_N(net291),
    .X(net297));
 sky130_fd_sc_hd__xnor2_4 c404 (.A(net292),
    .B(net294),
    .Y(net298));
 sky130_fd_sc_hd__xnor2_2 c405 (.A(net70),
    .B(net876),
    .Y(net299));
 sky130_fd_sc_hd__buf_1 c406 (.A(net664),
    .X(net300));
 sky130_fd_sc_hd__a31o_4 c407 (.A1(net70),
    .A2(net298),
    .A3(net297),
    .B1(net300),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 c408 (.A(net1006),
    .X(net909));
 sky130_fd_sc_hd__a21bo_1 c409 (.A1(net301),
    .A2(net300),
    .B1_N(net291),
    .X(net302));
 sky130_fd_sc_hd__a21bo_1 c410 (.A1(net297),
    .A2(net299),
    .B1_N(net291),
    .X(net303));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(net303),
    .A2(net193),
    .B1_N(net192),
    .X(net304));
 sky130_fd_sc_hd__a41o_1 c412 (.A1(net294),
    .A2(net909),
    .A3(net303),
    .A4(net945),
    .B1(net200),
    .X(net305));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net302),
    .A2(net293),
    .B1_N(net945),
    .X(net306));
 sky130_fd_sc_hd__a31o_1 c414 (.A1(net299),
    .A2(net297),
    .A3(net945),
    .B1(net909),
    .X(net307));
 sky130_fd_sc_hd__sdfsbp_2 c415 (.CLK(clknet_4_1_0_clk),
    .D(net307),
    .SCD(net305),
    .SCE(net302),
    .SET_B(net306),
    .Q(net309),
    .Q_N(net308));
 sky130_fd_sc_hd__a41o_1 c416 (.A1(net1007),
    .A2(net307),
    .A3(net302),
    .A4(net306),
    .B1(net297),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net306),
    .A1(net879),
    .A2(net295),
    .A3(net309),
    .S0(net307),
    .S1(net663),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 c418 (.A(net706),
    .X(net312));
 sky130_fd_sc_hd__buf_2 c419 (.A(net667),
    .X(net313));
 sky130_fd_sc_hd__xnor2_1 c420 (.A(net298),
    .B(net313),
    .Y(net314));
 sky130_fd_sc_hd__a21bo_4 c421 (.A1(net192),
    .A2(net313),
    .B1_N(net208),
    .X(net901));
 sky130_fd_sc_hd__xnor2_4 c422 (.A(net871),
    .B(net953),
    .Y(net315));
 sky130_fd_sc_hd__xnor2_1 c423 (.A(net852),
    .B(net315),
    .Y(net316));
 sky130_fd_sc_hd__clkbuf_1 c424 (.A(net1018),
    .X(net317));
 sky130_fd_sc_hd__xnor2_1 c425 (.A(net314),
    .B(net313),
    .Y(net318));
 sky130_fd_sc_hd__clkbuf_2 c426 (.A(net651),
    .X(net319));
 sky130_fd_sc_hd__xnor2_1 c427 (.A(net214),
    .B(net901),
    .Y(net320));
 sky130_fd_sc_hd__a21bo_2 c428 (.A1(net315),
    .A2(net220),
    .B1_N(net320),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 c429 (.A(net706),
    .X(net322));
 sky130_fd_sc_hd__a21bo_1 c430 (.A1(net92),
    .A2(net298),
    .B1_N(net319),
    .X(net323));
 sky130_fd_sc_hd__a31o_1 c431 (.A1(net322),
    .A2(net316),
    .A3(net312),
    .B1(net984),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c432 (.A0(net185),
    .A1(net313),
    .A2(net305),
    .A3(net321),
    .S0(net88),
    .S1(net901),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net320),
    .A1(net323),
    .A2(net92),
    .A3(net901),
    .S0(net185),
    .S1(clknet_1_0__leaf_net760),
    .X(net326));
 sky130_fd_sc_hd__a21bo_1 c434 (.A1(net326),
    .A2(net298),
    .B1_N(net321),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 c435 (.A(net705),
    .X(net328));
 sky130_fd_sc_hd__a41o_1 c436 (.A1(net316),
    .A2(net319),
    .A3(net312),
    .A4(net321),
    .B1(clknet_1_0__leaf_net760),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(net328),
    .A1(net937),
    .A2(clknet_1_0__leaf_net329),
    .A3(net324),
    .S0(clknet_1_0__leaf_net327),
    .S1(clknet_1_0__leaf_net760),
    .X(net330));
 sky130_fd_sc_hd__dlymetal6s2s_1 c438 (.A(net722),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net318),
    .A1(clknet_1_0__leaf_net329),
    .A2(net315),
    .A3(net92),
    .S0(net331),
    .S1(net322),
    .X(net332));
 sky130_fd_sc_hd__buf_1 c440 (.A(net723),
    .X(net333));
 sky130_fd_sc_hd__buf_1 c441 (.A(net723),
    .X(net334));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net333),
    .A2(net323),
    .B1_N(net861),
    .X(net335));
 sky130_fd_sc_hd__sdfsbp_1 c443 (.CLK(clknet_4_3_0_clk),
    .D(net313),
    .SCD(net333),
    .SCE(net119),
    .SET_B(net940),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__a21bo_1 c444 (.A1(net331),
    .A2(net337),
    .B1_N(net940),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net892),
    .A1(net239),
    .A2(net952),
    .A3(net231),
    .S0(net336),
    .S1(net940),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(net323),
    .A1(net331),
    .A2(net952),
    .A3(net315),
    .S0(net940),
    .S1(net750),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net338),
    .A1(net242),
    .A2(net941),
    .A3(net865),
    .S0(net319),
    .S1(net945),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net821),
    .A1(net334),
    .A2(net207),
    .A3(net340),
    .S0(net749),
    .S1(net761),
    .X(net342));
 sky130_fd_sc_hd__sdfbbn_1 c449 (.CLK_N(clknet_4_1_0_clk),
    .D(net340),
    .RESET_B(net319),
    .SCD(net315),
    .SCE(net861),
    .SET_B(net940),
    .Q(net344),
    .Q_N(net343));
 sky130_fd_sc_hd__sdfstp_1 c450 (.CLK(clknet_4_0_0_clk),
    .D(net309),
    .SCD(net340),
    .SCE(net940),
    .SET_B(net942),
    .Q(net345));
 sky130_fd_sc_hd__a21bo_2 c451 (.A1(net859),
    .A2(net343),
    .B1_N(net751),
    .X(net899));
 sky130_fd_sc_hd__mux4_2 c452 (.A0(net334),
    .A1(net331),
    .A2(net333),
    .A3(net235),
    .S0(net688),
    .S1(net764),
    .X(net346));
 sky130_fd_sc_hd__sdfbbp_1 c453 (.CLK(clknet_4_1_0_clk),
    .D(net324),
    .RESET_B(net1005),
    .SCD(net239),
    .SCE(net946),
    .SET_B(net940),
    .Q(net348),
    .Q_N(net347));
 sky130_fd_sc_hd__a21bo_1 c454 (.A1(net836),
    .A2(net324),
    .B1_N(net764),
    .X(net349));
 sky130_fd_sc_hd__buf_1 c455 (.A(net816),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net866),
    .A1(net231),
    .A2(net942),
    .A3(net346),
    .S0(net88),
    .S1(net236),
    .X(net351));
 sky130_fd_sc_hd__buf_2 c457 (.A(net1006),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net828),
    .A1(net197),
    .A2(net352),
    .A3(net865),
    .S0(net347),
    .S1(net765),
    .X(net353));
 sky130_fd_sc_hd__a21bo_1 c459 (.A1(net349),
    .A2(net899),
    .B1_N(net315),
    .X(net354));
 sky130_fd_sc_hd__a21bo_1 c460 (.A1(net334),
    .A2(net348),
    .B1_N(net345),
    .X(net355));
 sky130_fd_sc_hd__a21bo_1 c461 (.A1(net353),
    .A2(net355),
    .B1_N(net347),
    .X(net356));
 sky130_fd_sc_hd__a31o_1 c462 (.A1(net908),
    .A2(net112),
    .A3(net757),
    .B1(clknet_1_1__leaf_net760),
    .X(net357));
 sky130_fd_sc_hd__a31o_1 c463 (.A1(net299),
    .A2(net253),
    .A3(net352),
    .B1(net908),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 c464 (.A0(net253),
    .A1(net228),
    .A2(net133),
    .A3(net960),
    .S0(net867),
    .S1(net905),
    .X(net359));
 sky130_fd_sc_hd__buf_1 c465 (.A(net816),
    .X(net360));
 sky130_fd_sc_hd__a41o_1 c466 (.A1(net248),
    .A2(clknet_1_0__leaf_net262),
    .A3(net989),
    .A4(net139),
    .B1(net359),
    .X(net361));
 sky130_fd_sc_hd__a31o_1 c467 (.A1(net360),
    .A2(net346),
    .A3(net359),
    .B1(clknet_1_1__leaf_net357),
    .X(net362));
 sky130_fd_sc_hd__a31o_1 c468 (.A1(clknet_1_0__leaf_net357),
    .A2(net197),
    .A3(net941),
    .B1(net688),
    .X(net363));
 sky130_fd_sc_hd__a31o_1 c469 (.A1(net112),
    .A2(net854),
    .A3(clknet_1_1__leaf_net329),
    .B1(net229),
    .X(net364));
 sky130_fd_sc_hd__sdfbbn_1 c470 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_1__leaf_net262),
    .RESET_B(net88),
    .SCD(net990),
    .SCE(net133),
    .SET_B(net1012),
    .Q(net894),
    .Q_N(net365));
 sky130_fd_sc_hd__mux4_2 c471 (.A0(net140),
    .A1(net911),
    .A2(net133),
    .A3(net248),
    .S0(net112),
    .S1(net765),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net346),
    .A1(clknet_1_0__leaf_net363),
    .A2(net937),
    .A3(net867),
    .S0(net993),
    .S1(net749),
    .X(net367));
 sky130_fd_sc_hd__a31o_1 c473 (.A1(net854),
    .A2(net197),
    .A3(net952),
    .B1(net734),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net879),
    .A1(net253),
    .A2(clknet_1_0__leaf_net363),
    .A3(net993),
    .S0(net686),
    .S1(net734),
    .X(net369));
 sky130_fd_sc_hd__a31o_1 c475 (.A1(net236),
    .A2(clknet_1_0__leaf_net363),
    .A3(clknet_1_1__leaf_net357),
    .B1(net768),
    .X(net370));
 sky130_fd_sc_hd__sdfstp_1 c476 (.CLK(clknet_4_12_0_clk),
    .D(net368),
    .SCD(net346),
    .SCE(net360),
    .SET_B(net909),
    .Q(net371));
 sky130_fd_sc_hd__a41o_1 c477 (.A1(net352),
    .A2(net371),
    .A3(net718),
    .A4(net751),
    .B1(net766),
    .X(net372));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net876),
    .A2(net372),
    .A3(clknet_1_0__leaf_net363),
    .A4(net685),
    .B1(net768),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net228),
    .A1(clknet_1_0__leaf_net357),
    .A2(net372),
    .A3(net299),
    .S0(net346),
    .S1(net768),
    .X(net374));
 sky130_fd_sc_hd__a41o_1 c480 (.A1(net197),
    .A2(net974),
    .A3(net372),
    .A4(net371),
    .B1(net688),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net375),
    .A1(net348),
    .A2(net207),
    .A3(net909),
    .S0(net359),
    .S1(clknet_1_0__leaf_net363),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net371),
    .A1(net375),
    .A2(net372),
    .A3(clknet_1_0__leaf_net262),
    .S0(clknet_1_1__leaf_net760),
    .S1(net768),
    .X(net377));
 sky130_fd_sc_hd__mux4_2 c483 (.A0(net865),
    .A1(net371),
    .A2(net375),
    .A3(net939),
    .S0(net725),
    .S1(clknet_1_1__leaf_net759),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net263),
    .A1(net899),
    .A2(net876),
    .A3(net285),
    .S0(net880),
    .S1(net766),
    .X(net379));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(clknet_1_1__leaf_net329),
    .A1(clknet_1_0__leaf_net378),
    .A2(net829),
    .A3(net938),
    .S0(net893),
    .S1(net942),
    .X(net380));
 sky130_fd_sc_hd__sdfbbn_1 c486 (.CLK_N(clknet_4_14_0_clk),
    .D(net938),
    .RESET_B(net952),
    .SCD(net901),
    .SCE(net139),
    .SET_B(clknet_1_0__leaf_net378),
    .Q(net382),
    .Q_N(net381));
 sky130_fd_sc_hd__a41o_1 c487 (.A1(net278),
    .A2(net942),
    .A3(net897),
    .A4(net276),
    .B1(net765),
    .X(net383));
 sky130_fd_sc_hd__a41o_1 c488 (.A1(net383),
    .A2(net909),
    .A3(net867),
    .A4(net952),
    .B1(net962),
    .X(net384));
 sky130_fd_sc_hd__sdfbbp_1 c489 (.CLK(clknet_4_11_0_clk),
    .D(net276),
    .RESET_B(clknet_1_1__leaf_net378),
    .SCD(net365),
    .SCE(net860),
    .SET_B(net746),
    .Q(net907),
    .Q_N(net385));
 sky130_fd_sc_hd__sdfbbn_1 c490 (.CLK_N(clknet_4_14_0_clk),
    .D(net272),
    .RESET_B(clknet_1_0__leaf_net363),
    .SCD(net867),
    .SCE(net765),
    .SET_B(net888),
    .Q(net387),
    .Q_N(net386));
 sky130_fd_sc_hd__a41o_1 c491 (.A1(clknet_1_1__leaf_net256),
    .A2(net383),
    .A3(net920),
    .A4(net900),
    .B1(net769),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net901),
    .A1(net939),
    .A2(net285),
    .A3(net270),
    .S0(net666),
    .S1(net962),
    .X(net912));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(clknet_1_0__leaf_net283),
    .A1(net897),
    .A2(clknet_1_1__leaf_net378),
    .A3(net960),
    .S0(net263),
    .S1(net938),
    .X(net389));
 sky130_fd_sc_hd__a21bo_1 c494 (.A1(net168),
    .A2(net829),
    .B1_N(net270),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(clknet_1_1__leaf_net378),
    .A1(net991),
    .A2(net897),
    .A3(net942),
    .S0(net962),
    .S1(net770),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net897),
    .A1(net953),
    .A2(net861),
    .A3(net383),
    .S0(net768),
    .S1(net773),
    .X(net392));
 sky130_fd_sc_hd__a41o_1 c497 (.A1(net865),
    .A2(net938),
    .A3(net385),
    .A4(net757),
    .B1(net773),
    .X(net393));
 sky130_fd_sc_hd__a41o_2 c498 (.A1(net880),
    .A2(net29),
    .A3(net951),
    .A4(net962),
    .B1(net773),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net227),
    .A1(net387),
    .A2(net151),
    .A3(net897),
    .S0(clknet_1_1__leaf_net283),
    .S1(net772),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net160),
    .A1(net393),
    .A2(net394),
    .A3(net913),
    .S0(net962),
    .S1(net772),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(clknet_1_1__leaf_net251),
    .A1(net665),
    .A2(net962),
    .A3(net771),
    .S0(net773),
    .S1(net774),
    .X(net397));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(net390),
    .A1(net29),
    .A2(net167),
    .A3(net744),
    .S0(net927),
    .S1(net962),
    .X(net398));
 sky130_fd_sc_hd__a41o_1 c503 (.A1(net942),
    .A2(net398),
    .A3(net897),
    .A4(net898),
    .B1(net962),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net348),
    .A1(net398),
    .A2(net942),
    .A3(net115),
    .S0(net771),
    .S1(net772),
    .X(net400));
 sky130_fd_sc_hd__sdfbbn_2 c505 (.CLK_N(clknet_4_14_0_clk),
    .D(net398),
    .RESET_B(net993),
    .SCD(net1021),
    .SCE(net910),
    .SET_B(net772),
    .Q(net882),
    .Q_N(net401));
 sky130_fd_sc_hd__clkbuf_2 c528 (.A(net676),
    .X(net402));
 sky130_fd_sc_hd__a21bo_2 c529 (.A1(net194),
    .A2(net64),
    .B1_N(net402),
    .X(net403));
 sky130_fd_sc_hd__xnor2_4 c530 (.A(net67),
    .B(net301),
    .Y(net404));
 sky130_fd_sc_hd__mux4_2 c531 (.A0(net74),
    .A1(net291),
    .A2(net303),
    .A3(net194),
    .S0(net294),
    .S1(net663),
    .X(net405));
 sky130_fd_sc_hd__xnor2_1 c532 (.A(net818),
    .B(net404),
    .Y(net406));
 sky130_fd_sc_hd__xnor2_2 c533 (.A(net403),
    .B(net301),
    .Y(net407));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net187),
    .A1(net64),
    .A2(net404),
    .A3(net403),
    .S0(net402),
    .S1(net749),
    .X(net408));
 sky130_fd_sc_hd__xnor2_2 c535 (.A(net407),
    .B(net402),
    .Y(net409));
 sky130_fd_sc_hd__buf_1 c536 (.A(net676),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_4 c537 (.A(net705),
    .X(net411));
 sky130_fd_sc_hd__xnor2_4 c538 (.A(net404),
    .B(net411),
    .Y(net412));
 sky130_fd_sc_hd__xnor2_1 c539 (.A(net303),
    .B(net405),
    .Y(net413));
 sky130_fd_sc_hd__xnor2_1 c540 (.A(net410),
    .B(net664),
    .Y(net414));
 sky130_fd_sc_hd__xnor2_2 c541 (.A(net413),
    .B(net411),
    .Y(net415));
 sky130_fd_sc_hd__clkbuf_1 c542 (.A(net700),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 c543 (.A(net676),
    .X(net417));
 sky130_fd_sc_hd__xnor2_1 c544 (.A(net410),
    .B(net411),
    .Y(net418));
 sky130_fd_sc_hd__sdfstp_2 c545 (.CLK(clknet_4_4_0_clk),
    .D(net416),
    .SCD(net407),
    .SCE(net412),
    .SET_B(net405),
    .Q(net419));
 sky130_fd_sc_hd__buf_1 c546 (.A(net646),
    .X(net420));
 sky130_fd_sc_hd__xnor2_4 c547 (.A(net417),
    .B(net419),
    .Y(net421));
 sky130_fd_sc_hd__a31o_1 c548 (.A1(net419),
    .A2(net187),
    .A3(net421),
    .B1(net947),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net618),
    .A1(net419),
    .A2(net421),
    .A3(net422),
    .S0(net415),
    .S1(net879),
    .X(net423));
 sky130_fd_sc_hd__xnor2_4 c550 (.A(net309),
    .B(net312),
    .Y(net424));
 sky130_fd_sc_hd__buf_1 c551 (.A(net704),
    .X(net425));
 sky130_fd_sc_hd__xnor2_2 c552 (.A(net321),
    .B(net421),
    .Y(net426));
 sky130_fd_sc_hd__buf_1 c553 (.A(net815),
    .X(net427));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net420),
    .B(net403),
    .Y(net428));
 sky130_fd_sc_hd__dlymetal6s2s_1 c555 (.A(net638),
    .X(net429));
 sky130_fd_sc_hd__xnor2_1 c556 (.A(net427),
    .B(net414),
    .Y(net430));
 sky130_fd_sc_hd__xnor2_1 c557 (.A(net951),
    .B(net761),
    .Y(net431));
 sky130_fd_sc_hd__xnor2_1 c558 (.A(net425),
    .B(net74),
    .Y(net432));
 sky130_fd_sc_hd__clkbuf_4 c559 (.A(net815),
    .X(net886));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net220),
    .A1(net937),
    .A2(net886),
    .A3(net409),
    .S0(net411),
    .S1(net425),
    .X(net433));
 sky130_fd_sc_hd__a21bo_1 c561 (.A1(net428),
    .A2(net411),
    .B1_N(net414),
    .X(net434));
 sky130_fd_sc_hd__a21bo_1 c562 (.A1(net402),
    .A2(net220),
    .B1_N(clknet_1_0__leaf_net760),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 c563 (.A(net722),
    .X(net436));
 sky130_fd_sc_hd__a21bo_1 c564 (.A1(net434),
    .A2(net427),
    .B1_N(net776),
    .X(net437));
 sky130_fd_sc_hd__buf_2 c565 (.A(net638),
    .X(net438));
 sky130_fd_sc_hd__a31o_1 c566 (.A1(net436),
    .A2(net886),
    .A3(net437),
    .B1(net776),
    .X(net439));
 sky130_fd_sc_hd__xnor2_2 c567 (.A(net439),
    .B(net420),
    .Y(net440));
 sky130_fd_sc_hd__buf_1 c568 (.A(net650),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net432),
    .A1(net436),
    .A2(net438),
    .A3(net937),
    .S0(net886),
    .S1(net1010),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net414),
    .A1(net439),
    .A2(net434),
    .A3(net312),
    .S0(net440),
    .S1(net776),
    .X(net443));
 sky130_fd_sc_hd__sdfbbp_1 c571 (.CLK(clknet_4_4_0_clk),
    .D(net431),
    .RESET_B(net440),
    .SCD(net425),
    .SCE(net441),
    .SET_B(net1004),
    .Q(net445),
    .Q_N(net444));
 sky130_fd_sc_hd__buf_2 c572 (.A(net814),
    .X(net446));
 sky130_fd_sc_hd__a21bo_1 c573 (.A1(net403),
    .A2(net446),
    .B1_N(net354),
    .X(net447));
 sky130_fd_sc_hd__a41o_1 c574 (.A1(net441),
    .A2(net829),
    .A3(net405),
    .A4(net984),
    .B1(net776),
    .X(net448));
 sky130_fd_sc_hd__sdfbbn_1 c575 (.CLK_N(clknet_4_1_0_clk),
    .D(net447),
    .RESET_B(net947),
    .SCD(net677),
    .SCE(clknet_1_0__leaf_net760),
    .SET_B(net775),
    .Q(net450),
    .Q_N(net449));
 sky130_fd_sc_hd__a41o_2 c576 (.A1(net231),
    .A2(net860),
    .A3(net356),
    .A4(net308),
    .B1(net756),
    .X(net451));
 sky130_fd_sc_hd__a41o_1 c577 (.A1(net354),
    .A2(net886),
    .A3(net239),
    .A4(net231),
    .B1(net677),
    .X(net452));
 sky130_fd_sc_hd__buf_1 c578 (.A(net814),
    .X(net453));
 sky130_fd_sc_hd__a41o_1 c579 (.A1(net241),
    .A2(net344),
    .A3(net441),
    .A4(net750),
    .B1(net766),
    .X(net454));
 sky130_fd_sc_hd__sedfxbp_1 c580 (.CLK(clknet_4_4_0_clk),
    .D(net447),
    .DE(net450),
    .SCD(net207),
    .SCE(net424),
    .Q(net456),
    .Q_N(net455));
 sky130_fd_sc_hd__a41o_2 c581 (.A1(net456),
    .A2(net405),
    .A3(net449),
    .A4(net453),
    .B1(net756),
    .X(net877));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net441),
    .A1(net886),
    .A2(net350),
    .A3(clknet_1_0__leaf_net760),
    .S0(net762),
    .S1(net775),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net448),
    .A1(clknet_1_1__leaf_net457),
    .A2(net953),
    .A3(net446),
    .S0(net750),
    .S1(net775),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net829),
    .A1(net409),
    .A2(net447),
    .A3(net231),
    .S0(net729),
    .S1(net775),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net355),
    .A1(clknet_1_0__leaf_net458),
    .A2(net405),
    .A3(net877),
    .S0(net446),
    .S1(net242),
    .X(net460));
 sky130_fd_sc_hd__sdfbbn_1 c586 (.CLK_N(clknet_4_3_0_clk),
    .D(net337),
    .RESET_B(clknet_1_0__leaf_net458),
    .SCD(net1025),
    .SCE(net761),
    .SET_B(clknet_1_0__leaf_net778),
    .Q(net462),
    .Q_N(net461));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_0__leaf_net457),
    .A1(net231),
    .A2(clknet_1_1__leaf_net458),
    .A3(net447),
    .S0(net455),
    .S1(clknet_1_1__leaf_net778),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net344),
    .A1(net877),
    .A2(clknet_1_1__leaf_net458),
    .A3(net451),
    .S0(clknet_1_0__leaf_net777),
    .S1(clknet_1_0__leaf_net779),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net409),
    .A1(clknet_1_1__leaf_net458),
    .A2(clknet_1_1__leaf_net435),
    .A3(net355),
    .S0(net953),
    .S1(clknet_1_1__leaf_net779),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net461),
    .A1(net945),
    .A2(clknet_1_0__leaf_net458),
    .A3(net756),
    .S0(clknet_1_1__leaf_net777),
    .S1(net780),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net453),
    .A1(net438),
    .A2(net451),
    .A3(clknet_1_1__leaf_net458),
    .S0(net446),
    .S1(net424),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net447),
    .A1(net694),
    .A2(net766),
    .A3(net781),
    .S0(net782),
    .S1(net784),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net239),
    .A1(net462),
    .A2(net877),
    .A3(clknet_1_0__leaf_net458),
    .S0(clknet_1_0__leaf_net703),
    .S1(net784),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net105),
    .A1(net877),
    .A2(net948),
    .A3(net82),
    .S0(net953),
    .S1(net767),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(clknet_1_0__leaf_net357),
    .A1(net260),
    .A2(net146),
    .A3(net133),
    .S0(net940),
    .S1(net964),
    .X(net471));
 sky130_fd_sc_hd__sedfxbp_1 c596 (.CLK(clknet_4_12_0_clk),
    .D(net207),
    .DE(net899),
    .SCD(net259),
    .SCE(net993),
    .Q(net473),
    .Q_N(net472));
 sky130_fd_sc_hd__sedfxtp_1 c597 (.CLK(clknet_4_3_0_clk),
    .D(net260),
    .DE(net105),
    .SCD(net824),
    .SCE(net775),
    .Q(net474));
 sky130_fd_sc_hd__mux4_2 c598 (.A0(net473),
    .A1(net125),
    .A2(net939),
    .A3(net958),
    .S0(net259),
    .S1(net767),
    .X(net475));
 sky130_fd_sc_hd__a31o_1 c599 (.A1(net474),
    .A2(clknet_1_1__leaf_net357),
    .A3(net259),
    .B1(net775),
    .X(net476));
 sky130_fd_sc_hd__a41o_2 c600 (.A1(net372),
    .A2(net125),
    .A3(net939),
    .A4(net964),
    .B1(net775),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net476),
    .A1(net879),
    .A2(net865),
    .A3(net940),
    .S0(net749),
    .S1(net776),
    .X(net478));
 sky130_fd_sc_hd__a31o_1 c602 (.A1(net429),
    .A2(net941),
    .A3(clknet_1_0__leaf_net759),
    .B1(clknet_1_1__leaf_net760),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net350),
    .A1(clknet_1_1__leaf_net479),
    .A2(clknet_1_0__leaf_net478),
    .A3(net474),
    .S0(net984),
    .S1(net776),
    .X(net480));
 sky130_fd_sc_hd__sdfbbp_1 c604 (.CLK(clknet_4_6_0_clk),
    .D(net444),
    .RESET_B(net936),
    .SCD(net957),
    .SCE(net689),
    .SET_B(net1001),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net123),
    .A1(net304),
    .A2(net936),
    .A3(clknet_1_0__leaf_net478),
    .S0(net964),
    .S1(net775),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net147),
    .A1(clknet_1_0__leaf_net478),
    .A2(net372),
    .A3(net123),
    .S0(net936),
    .S1(net946),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net450),
    .A1(clknet_1_0__leaf_net471),
    .A2(net936),
    .A3(net993),
    .S0(net940),
    .S1(net123),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net424),
    .A1(net260),
    .A2(net939),
    .A3(net359),
    .S0(net475),
    .S1(net1024),
    .X(net486));
 sky130_fd_sc_hd__sedfxtp_4 c609 (.CLK(clknet_4_12_0_clk),
    .D(net125),
    .DE(net936),
    .SCD(net786),
    .SCE(net1026),
    .Q(net883));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net260),
    .A1(net948),
    .A2(net207),
    .A3(clknet_1_1__leaf_net471),
    .S0(clknet_1_1__leaf_net703),
    .S1(net786),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net482),
    .A1(net936),
    .A2(net472),
    .A3(net207),
    .S0(net788),
    .S1(net790),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net909),
    .A1(net883),
    .A2(net449),
    .A3(net775),
    .S0(net790),
    .S1(net792),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net883),
    .A1(net936),
    .A2(net957),
    .A3(net689),
    .S0(net963),
    .S1(net1022),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net489),
    .A1(net481),
    .A2(net776),
    .A3(net789),
    .S0(net791),
    .S1(net793),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net242),
    .A1(net491),
    .A2(clknet_1_0__leaf_net479),
    .A3(net424),
    .S0(net791),
    .S1(net793),
    .X(net492));
 sky130_fd_sc_hd__sedfxtp_1 c616 (.CLK(clknet_4_14_0_clk),
    .D(net429),
    .DE(net359),
    .SCD(net1019),
    .SCE(net794),
    .Q(net493));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(clknet_1_1__leaf_net478),
    .A1(net445),
    .A2(net879),
    .A3(net909),
    .S0(net352),
    .S1(net151),
    .X(net494));
 sky130_fd_sc_hd__a31o_1 c618 (.A1(net151),
    .A2(net882),
    .A3(net957),
    .B1(net694),
    .X(net933));
 sky130_fd_sc_hd__sdfrbp_1 c619 (.CLK(clknet_4_15_0_clk),
    .D(net270),
    .RESET_B(net359),
    .SCD(net766),
    .SCE(net787),
    .Q(net496),
    .Q_N(net495));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net833),
    .A1(net830),
    .A2(net845),
    .A3(net3),
    .S0(net868),
    .S1(net854),
    .X(net0));
 sky130_fd_sc_hd__sdfbbn_1 c620 (.CLK_N(clknet_4_12_0_clk),
    .D(clknet_1_1__leaf_net397),
    .RESET_B(net880),
    .SCD(net887),
    .SCE(net444),
    .SET_B(net899),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net270),
    .A1(net379),
    .A2(net401),
    .A3(net886),
    .S0(clknet_1_1__leaf_net759),
    .S1(net794),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net958),
    .A1(clknet_1_0__leaf_net889),
    .A2(net270),
    .A3(net935),
    .S0(net787),
    .S1(net794),
    .X(net499));
 sky130_fd_sc_hd__a31o_1 c623 (.A1(net88),
    .A2(net82),
    .A3(net497),
    .B1(net958),
    .X(net890));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(clknet_1_0__leaf_net363),
    .A1(net495),
    .A2(net270),
    .A3(net951),
    .S0(clknet_1_1__leaf_net478),
    .X(net500));
 sky130_fd_sc_hd__a41o_1 c625 (.A1(net951),
    .A2(net886),
    .A3(net270),
    .A4(net962),
    .B1(net794),
    .X(net501));
 sky130_fd_sc_hd__a41o_1 c626 (.A1(net860),
    .A2(net401),
    .A3(net690),
    .A4(net694),
    .B1(net794),
    .X(net502));
 sky130_fd_sc_hd__a31o_1 c627 (.A1(net496),
    .A2(net876),
    .A3(net270),
    .B1(net774),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net359),
    .A1(net882),
    .A2(net493),
    .A3(net501),
    .S0(net285),
    .S1(net1023),
    .X(net504));
 sky130_fd_sc_hd__a41o_1 c629 (.A1(net977),
    .A2(net379),
    .A3(net493),
    .A4(net861),
    .B1(net860),
    .X(net505));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net870),
    .A1(net873),
    .A2(net867),
    .A3(net0),
    .S0(net855),
    .S1(net868),
    .X(net1));
 sky130_fd_sc_hd__sdfbbn_2 c630 (.CLK_N(clknet_4_14_0_clk),
    .D(net1011),
    .RESET_B(net493),
    .SCD(clknet_1_0__leaf_net889),
    .SCE(net501),
    .SET_B(net359),
    .Q(net507),
    .Q_N(net506));
 sky130_fd_sc_hd__a41o_1 c631 (.A1(net133),
    .A2(net505),
    .A3(net501),
    .A4(net506),
    .B1(net795),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net503),
    .A1(net507),
    .A2(net501),
    .A3(net401),
    .S0(net505),
    .S1(net769),
    .X(net509));
 sky130_fd_sc_hd__a31o_1 c633 (.A1(net352),
    .A2(net502),
    .A3(net507),
    .B1(net962),
    .X(net510));
 sky130_fd_sc_hd__a31o_1 c634 (.A1(net498),
    .A2(net507),
    .A3(net794),
    .B1(net795),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net511),
    .A1(net502),
    .A2(net381),
    .A3(net506),
    .S0(net745),
    .S1(clknet_1_1__leaf_net759),
    .X(net512));
 sky130_fd_sc_hd__a31o_1 c636 (.A1(net510),
    .A2(net501),
    .A3(net882),
    .B1(net511),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net860),
    .A1(net512),
    .A2(net507),
    .A3(net513),
    .S0(clknet_1_0__leaf_net397),
    .S1(net795),
    .X(net514));
 sky130_fd_sc_hd__mux4_1 c64 (.A0(net856),
    .A1(net876),
    .A2(net868),
    .A3(net866),
    .S0(net830),
    .S1(net865),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c65 (.A0(net871),
    .A1(net847),
    .A2(net840),
    .A3(net835),
    .S0(net845),
    .S1(net823),
    .X(net3));
 sky130_fd_sc_hd__xnor2_2 c66 (.A(net860),
    .B(net834),
    .Y(net4));
 sky130_fd_sc_hd__clkbuf_2 c660 (.A(net700),
    .X(net515));
 sky130_fd_sc_hd__a21bo_1 c661 (.A1(net301),
    .A2(net422),
    .B1_N(clknet_1_0__leaf_net759),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_1 c662 (.A(net682),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_4 c663 (.A(net682),
    .X(net518));
 sky130_fd_sc_hd__buf_4 c664 (.A(net719),
    .X(net519));
 sky130_fd_sc_hd__buf_1 c665 (.A(net700),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_2 c666 (.A(net646),
    .X(net521));
 sky130_fd_sc_hd__mux4_2 c667 (.A0(net961),
    .A1(net404),
    .A2(net301),
    .A3(net292),
    .S0(net518),
    .S1(net519),
    .X(net522));
 sky130_fd_sc_hd__xnor2_1 c668 (.A(net517),
    .B(clknet_1_0__leaf_net759),
    .Y(net523));
 sky130_fd_sc_hd__sdfrbp_1 c669 (.CLK(clknet_4_5_0_clk),
    .D(net294),
    .RESET_B(net522),
    .SCD(net518),
    .SCE(net520),
    .Q(net525),
    .Q_N(net524));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net867),
    .B(net968),
    .Y(net5));
 sky130_fd_sc_hd__a31o_1 c670 (.A1(net518),
    .A2(net200),
    .A3(net515),
    .B1(net519),
    .X(net526));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net945),
    .A1(net522),
    .A2(net406),
    .A3(net519),
    .S0(net291),
    .S1(net961),
    .X(net527));
 sky130_fd_sc_hd__xnor2_1 c672 (.A(net518),
    .B(net683),
    .Y(net528));
 sky130_fd_sc_hd__buf_1 c673 (.A(net720),
    .X(net529));
 sky130_fd_sc_hd__xnor2_2 c674 (.A(net1020),
    .B(net683),
    .Y(net530));
 sky130_fd_sc_hd__xnor2_1 c675 (.A(net530),
    .B(net968),
    .Y(net531));
 sky130_fd_sc_hd__xnor2_2 c676 (.A(net529),
    .B(net519),
    .Y(net532));
 sky130_fd_sc_hd__buf_1 c677 (.A(net719),
    .X(net533));
 sky130_fd_sc_hd__xnor2_1 c678 (.A(net528),
    .B(net521),
    .Y(net534));
 sky130_fd_sc_hd__buf_1 c679 (.A(net676),
    .X(net535));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net835),
    .B(net5),
    .Y(net6));
 sky130_fd_sc_hd__buf_1 c680 (.A(net720),
    .X(net536));
 sky130_fd_sc_hd__a31o_1 c681 (.A1(net533),
    .A2(net530),
    .A3(net532),
    .B1(net518),
    .X(net537));
 sky130_fd_sc_hd__xnor2_1 c682 (.A(net535),
    .B(clknet_1_0__leaf_net435),
    .Y(net538));
 sky130_fd_sc_hd__a21bo_1 c683 (.A1(net200),
    .A2(net438),
    .B1_N(net530),
    .X(net539));
 sky130_fd_sc_hd__a31o_1 c684 (.A1(net421),
    .A2(clknet_1_0__leaf_net523),
    .A3(net968),
    .B1(net438),
    .X(net540));
 sky130_fd_sc_hd__a41o_1 c685 (.A1(net536),
    .A2(clknet_1_0__leaf_net435),
    .A3(net518),
    .A4(clknet_1_0__leaf_net540),
    .B1(clknet_1_0__leaf_net759),
    .X(net541));
 sky130_fd_sc_hd__a21bo_1 c686 (.A1(clknet_1_0__leaf_net540),
    .A2(net312),
    .B1_N(net421),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 c687 (.A(net704),
    .X(net543));
 sky130_fd_sc_hd__a21bo_1 c688 (.A1(net291),
    .A2(net537),
    .B1_N(net531),
    .X(net544));
 sky130_fd_sc_hd__a21bo_1 c689 (.A1(net312),
    .A2(clknet_1_0__leaf_net435),
    .B1_N(net762),
    .X(net545));
 sky130_fd_sc_hd__xnor2_1 c69 (.A(net2),
    .B(net4),
    .Y(net7));
 sky130_fd_sc_hd__a21bo_1 c690 (.A1(net541),
    .A2(clknet_1_0__leaf_net542),
    .B1_N(clknet_1_0__leaf_net435),
    .X(net546));
 sky130_fd_sc_hd__a21bo_1 c691 (.A1(net537),
    .A2(net945),
    .B1_N(net525),
    .X(net547));
 sky130_fd_sc_hd__a21bo_2 c692 (.A1(net543),
    .A2(net532),
    .B1_N(net530),
    .X(net548));
 sky130_fd_sc_hd__a41o_1 c693 (.A1(clknet_1_0__leaf_net542),
    .A2(net200),
    .A3(net537),
    .A4(clknet_1_1__leaf_net540),
    .B1(net532),
    .X(net549));
 sky130_fd_sc_hd__a31o_1 c694 (.A1(net545),
    .A2(clknet_1_0__leaf_net540),
    .A3(net544),
    .B1(net547),
    .X(net550));
 sky130_fd_sc_hd__a41o_1 c695 (.A1(net549),
    .A2(net519),
    .A3(clknet_1_1__leaf_net542),
    .A4(net522),
    .B1(net548),
    .X(net551));
 sky130_fd_sc_hd__sdfbbp_1 c696 (.CLK(clknet_4_5_0_clk),
    .D(net1020),
    .RESET_B(net548),
    .SCD(clknet_1_0__leaf_net435),
    .SCE(net519),
    .SET_B(clknet_1_1__leaf_net546),
    .Q(net553),
    .Q_N(net552));
 sky130_fd_sc_hd__a41o_1 c697 (.A1(net520),
    .A2(net438),
    .A3(net532),
    .A4(clknet_1_1__leaf_net542),
    .B1(net965),
    .X(net554));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(net530),
    .A2(clknet_1_1__leaf_net540),
    .A3(net312),
    .B1(net965),
    .X(net555));
 sky130_fd_sc_hd__a41o_1 c699 (.A1(net412),
    .A2(clknet_1_1__leaf_net546),
    .A3(net966),
    .A4(net548),
    .B1(net953),
    .X(net556));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net857),
    .B(net6),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net548),
    .A1(clknet_1_1__leaf_net554),
    .A2(clknet_1_1__leaf_net542),
    .A3(net966),
    .S0(net674),
    .S1(net762),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net540),
    .A1(clknet_1_1__leaf_net546),
    .A2(clknet_1_0__leaf_net557),
    .A3(net521),
    .S0(clknet_1_0__leaf_net554),
    .S1(net548),
    .X(net558));
 sky130_fd_sc_hd__a41o_1 c702 (.A1(clknet_1_0__leaf_net557),
    .A2(clknet_1_0__leaf_net554),
    .A3(net438),
    .A4(net548),
    .B1(net965),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net548),
    .A1(clknet_1_1__leaf_net557),
    .A2(net412),
    .A3(net524),
    .S0(clknet_1_0__leaf_net559),
    .S1(net719),
    .X(net560));
 sky130_fd_sc_hd__sdfbbn_1 c704 (.CLK_N(clknet_4_4_0_clk),
    .D(net235),
    .RESET_B(net446),
    .SCD(net119),
    .SCE(net965),
    .SET_B(net941),
    .Q(net562),
    .Q_N(net561));
 sky130_fd_sc_hd__a41o_1 c705 (.A1(clknet_1_0__leaf_net559),
    .A2(net451),
    .A3(net861),
    .A4(net963),
    .B1(clknet_1_0__leaf_net796),
    .X(net563));
 sky130_fd_sc_hd__mux4_2 c706 (.A0(net562),
    .A1(net984),
    .A2(net405),
    .A3(net544),
    .S0(net536),
    .S1(net963),
    .X(net564));
 sky130_fd_sc_hd__a41o_1 c707 (.A1(net876),
    .A2(net451),
    .A3(net966),
    .A4(net82),
    .B1(clknet_1_0__leaf_net796),
    .X(net565));
 sky130_fd_sc_hd__a41o_1 c708 (.A1(clknet_1_0__leaf_net565),
    .A2(net515),
    .A3(net562),
    .A4(net521),
    .B1(net966),
    .X(net566));
 sky130_fd_sc_hd__sdfbbn_1 c709 (.CLK_N(clknet_4_5_0_clk),
    .D(clknet_1_0__leaf_net546),
    .RESET_B(net521),
    .SCD(net966),
    .SCE(net235),
    .SET_B(net201),
    .Q(net568),
    .Q_N(net567));
 sky130_fd_sc_hd__xnor2_2 c71 (.A(net8),
    .B(net829),
    .Y(net9));
 sky130_fd_sc_hd__sdfbbp_1 c710 (.CLK(clknet_4_6_0_clk),
    .D(net448),
    .RESET_B(net438),
    .SCD(net235),
    .SCE(net88),
    .SET_B(clknet_1_1__leaf_net565),
    .Q(net570),
    .Q_N(net569));
 sky130_fd_sc_hd__a41o_1 c711 (.A1(net547),
    .A2(net567),
    .A3(net861),
    .A4(net966),
    .B1(net958),
    .X(net571));
 sky130_fd_sc_hd__sdfbbn_1 c712 (.CLK_N(clknet_4_7_0_clk),
    .D(net548),
    .RESET_B(net1003),
    .SCD(clknet_1_0__leaf_net563),
    .SCE(net451),
    .SET_B(net547),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__a41o_1 c713 (.A1(net521),
    .A2(net571),
    .A3(net223),
    .A4(net965),
    .B1(net783),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net536),
    .A1(net568),
    .A2(clknet_1_0__leaf_net546),
    .A3(net515),
    .S0(net82),
    .S1(net965),
    .X(net575));
 sky130_fd_sc_hd__a41o_1 c715 (.A1(net571),
    .A2(net573),
    .A3(net521),
    .A4(clknet_1_0__leaf_net538),
    .B1(net947),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net405),
    .A1(clknet_1_0__leaf_net546),
    .A2(net571),
    .A3(net958),
    .S0(net522),
    .S1(clknet_1_0__leaf_net797),
    .X(net577));
 sky130_fd_sc_hd__sdfrtn_1 c717 (.CLK_N(clknet_4_6_0_clk),
    .D(net119),
    .RESET_B(net998),
    .SCD(net965),
    .SCE(clknet_1_0__leaf_net703),
    .Q(net578));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net550),
    .A1(net946),
    .A2(net945),
    .A3(net966),
    .S0(clknet_1_0__leaf_net565),
    .S1(clknet_1_1__leaf_net797),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_1__leaf_net523),
    .A1(net438),
    .A2(net519),
    .A3(net762),
    .S0(clknet_1_0__leaf_net796),
    .S1(net800),
    .X(net580));
 sky130_fd_sc_hd__xnor2_1 c72 (.A(net864),
    .B(net870),
    .Y(net10));
 sky130_fd_sc_hd__a41o_1 c720 (.A1(net564),
    .A2(net515),
    .A3(net721),
    .A4(net785),
    .B1(net800),
    .X(net581));
 sky130_fd_sc_hd__a41o_1 c721 (.A1(net531),
    .A2(net451),
    .A3(net573),
    .A4(net548),
    .B1(net966),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net515),
    .A1(net580),
    .A2(net582),
    .A3(net119),
    .S0(net965),
    .S1(net581),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net581),
    .A1(net515),
    .A2(net544),
    .A3(clknet_1_0__leaf_net538),
    .S0(net673),
    .S1(clknet_1_0__leaf_net798),
    .X(net584));
 sky130_fd_sc_hd__sdfbbn_1 c724 (.CLK_N(clknet_4_7_0_clk),
    .D(net539),
    .RESET_B(net582),
    .SCD(clknet_1_1__leaf_net559),
    .SCE(net965),
    .SET_B(net804),
    .Q(net586),
    .Q_N(net585));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net555),
    .A1(net582),
    .A2(clknet_1_0__leaf_net563),
    .A3(net572),
    .S0(net561),
    .S1(net803),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(clknet_1_1__leaf_net563),
    .A1(net941),
    .A2(net936),
    .A3(clknet_1_1__leaf_net435),
    .S0(clknet_1_1__leaf_net363),
    .S1(clknet_1_1__leaf_net796),
    .X(net588));
 sky130_fd_sc_hd__a41o_1 c727 (.A1(net223),
    .A2(clknet_1_1__leaf_net563),
    .A3(clknet_1_1__leaf_net435),
    .A4(net793),
    .B1(net802),
    .X(net589));
 sky130_fd_sc_hd__a41o_1 c728 (.A1(net827),
    .A2(net586),
    .A3(net829),
    .A4(net936),
    .B1(net861),
    .X(net590));
 sky130_fd_sc_hd__a41o_1 c729 (.A1(net569),
    .A2(net729),
    .A3(net767),
    .A4(clknet_1_1__leaf_net796),
    .B1(net805),
    .X(net591));
 sky130_fd_sc_hd__xnor2_4 c73 (.A(net979),
    .B(net872),
    .Y(net11));
 sky130_fd_sc_hd__a41o_1 c730 (.A1(net578),
    .A2(net82),
    .A3(clknet_1_0__leaf_net591),
    .A4(net741),
    .B1(net799),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net936),
    .A1(clknet_1_1__leaf_net363),
    .A2(net519),
    .A3(clknet_1_1__leaf_net591),
    .S0(net223),
    .S1(net801),
    .X(net593));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net966),
    .A1(clknet_1_0__leaf_net591),
    .A2(net941),
    .A3(net948),
    .S0(net741),
    .S1(net807),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(clknet_1_1__leaf_net435),
    .A1(net592),
    .A2(net865),
    .A3(net477),
    .S0(net522),
    .S1(net805),
    .X(net595));
 sky130_fd_sc_hd__sdfbbp_1 c734 (.CLK(clknet_4_7_0_clk),
    .D(net957),
    .RESET_B(net522),
    .SCD(net1008),
    .SCE(clknet_1_1__leaf_net798),
    .SET_B(net807),
    .Q(net596));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net941),
    .A1(net570),
    .A2(net585),
    .A3(net946),
    .S0(net477),
    .S1(clknet_1_0__leaf_net798),
    .X(net597));
 sky130_fd_sc_hd__a31o_2 c736 (.A1(net966),
    .A2(net564),
    .A3(net729),
    .B1(net807),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net223),
    .A1(clknet_1_1__leaf_net563),
    .A2(net965),
    .A3(net709),
    .S0(net767),
    .S1(net807),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(clknet_1_1__leaf_net591),
    .A1(net941),
    .A2(net552),
    .A3(net710),
    .S0(net963),
    .S1(net806),
    .X(net600));
 sky130_fd_sc_hd__sdfbbn_1 c739 (.CLK_N(clknet_4_13_0_clk),
    .D(net600),
    .RESET_B(net553),
    .SCD(clknet_1_1__leaf_net363),
    .SCE(net689),
    .SET_B(clknet_1_1__leaf_net759),
    .Q(net601));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net996),
    .B(net870),
    .Y(net12));
 sky130_fd_sc_hd__sdfbbn_1 c740 (.CLK_N(clknet_4_7_0_clk),
    .D(net594),
    .RESET_B(net477),
    .SCD(net598),
    .SCE(net721),
    .SET_B(clknet_1_0__leaf_net796),
    .Q(net603),
    .Q_N(net602));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(net603),
    .A1(net596),
    .A2(net578),
    .A3(net564),
    .S0(clknet_1_1__leaf_net591),
    .S1(net807),
    .X(net604));
 sky130_fd_sc_hd__sdfbbp_1 c742 (.CLK(clknet_4_7_0_clk),
    .D(net518),
    .RESET_B(net603),
    .SCD(net598),
    .SCE(net793),
    .SET_B(net802),
    .Q(net605));
 sky130_fd_sc_hd__sdfbbn_1 c743 (.CLK_N(clknet_4_6_0_clk),
    .D(net1002),
    .RESET_B(clknet_1_0__leaf_net591),
    .SCD(net518),
    .SCE(net602),
    .SET_B(net598),
    .Q(net607),
    .Q_N(net606));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(clknet_1_1__leaf_net538),
    .A1(net598),
    .A2(net606),
    .A3(net793),
    .S0(clknet_1_1__leaf_net796),
    .S1(net799),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net604),
    .A1(net519),
    .A2(net603),
    .A3(net606),
    .S0(net713),
    .S1(net806),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net544),
    .A1(net605),
    .A2(net607),
    .A3(net602),
    .S0(clknet_1_1__leaf_net363),
    .S1(net808),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net607),
    .A1(net957),
    .A2(net712),
    .A3(net719),
    .S0(clknet_1_1__leaf_net796),
    .S1(net808),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net573),
    .A1(net522),
    .A2(net865),
    .A3(net394),
    .S0(net788),
    .S1(net808),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net519),
    .A1(net285),
    .A2(net475),
    .A3(net445),
    .S0(net82),
    .S1(net394),
    .X(net613));
 sky130_fd_sc_hd__a31o_4 c75 (.A1(net8),
    .A2(net10),
    .A3(net823),
    .B1(net845),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net446),
    .A1(net444),
    .A2(net394),
    .A3(net506),
    .S0(net729),
    .S1(net1013),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net475),
    .A1(net948),
    .A2(net860),
    .A3(net606),
    .S0(net732),
    .S1(net745),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net445),
    .A1(net394),
    .A2(net598),
    .A3(net506),
    .S0(clknet_1_1__leaf_net363),
    .S1(net963),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net867),
    .A1(net507),
    .A2(net732),
    .A3(net805),
    .S0(net808),
    .S1(net809),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net598),
    .A1(net88),
    .A2(net475),
    .A3(net564),
    .S1(net810),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net522),
    .A1(net946),
    .A2(net513),
    .A3(net607),
    .S0(net475),
    .S1(net598),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net564),
    .A1(net507),
    .A2(net445),
    .A3(net788),
    .S0(net999),
    .S1(net1030),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net572),
    .A1(net394),
    .A2(clknet_1_1__leaf_net703),
    .A3(net785),
    .S0(net810),
    .S1(net813),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net617),
    .A1(net611),
    .A2(net606),
    .A3(net800),
    .S0(net808),
    .S1(net813),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net506),
    .A1(net607),
    .A2(net695),
    .A3(net788),
    .S0(net808),
    .S1(net999),
    .X(net623));
 sky130_fd_sc_hd__a21bo_4 c76 (.A1(net9),
    .A2(net7),
    .B1_N(net954),
    .X(net14));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net957),
    .A1(net620),
    .A2(net861),
    .A3(net623),
    .S0(net1027),
    .S1(net999),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net622),
    .A1(net623),
    .A2(net598),
    .A3(net710),
    .S0(net718),
    .S1(net733),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net607),
    .A1(net394),
    .A2(net623),
    .A3(net709),
    .S0(net805),
    .S1(net812),
    .X(net626));
 sky130_fd_sc_hd__a31o_4 c77 (.A1(net870),
    .A2(net14),
    .A3(net6),
    .B1(net954),
    .X(net15));
 sky130_fd_sc_hd__a41o_1 c78 (.A1(net15),
    .A2(net856),
    .A3(net6),
    .A4(net867),
    .B1(net954),
    .X(net16));
 sky130_fd_sc_hd__a21bo_4 c79 (.A1(net851),
    .A2(net15),
    .B1_N(net954),
    .X(net17));
 sky130_fd_sc_hd__a21bo_1 c80 (.A1(net11),
    .A2(net17),
    .B1_N(net954),
    .X(net18));
 sky130_fd_sc_hd__mux4_1 c81 (.A0(net823),
    .A1(net9),
    .A2(net862),
    .A3(net954),
    .S0(net4),
    .S1(net14),
    .X(net19));
 sky130_fd_sc_hd__a31o_4 c82 (.A1(net16),
    .A2(net17),
    .A3(net12),
    .B1(net995),
    .X(net20));
 sky130_fd_sc_hd__a41o_4 c83 (.A1(net20),
    .A2(net19),
    .A3(net15),
    .A4(net18),
    .B1(net995),
    .X(net21));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net21),
    .A1(net20),
    .A2(net14),
    .A3(net856),
    .S0(net6),
    .S1(net995),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c85 (.A0(net15),
    .A1(net18),
    .A2(net22),
    .A3(net20),
    .S0(net869),
    .S1(net955),
    .X(net23));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net16),
    .A1(net854),
    .A2(net10),
    .A3(net22),
    .S0(net23),
    .S1(net20),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net4),
    .A1(net24),
    .A2(net21),
    .A3(net22),
    .S0(net955),
    .S1(net23),
    .X(net911));
 sky130_fd_sc_hd__xnor2_4 c88 (.A(net824),
    .B(net986),
    .Y(net25));
 sky130_fd_sc_hd__xnor2_1 c89 (.A(net9),
    .B(net983),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net834),
    .B(net873),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_2 c91 (.A(net21),
    .B(net861),
    .Y(net28));
 sky130_fd_sc_hd__a31o_1 c92 (.A1(net28),
    .A2(net944),
    .A3(net847),
    .B1(net856),
    .X(net29));
 sky130_fd_sc_hd__xnor2_1 c93 (.A(net25),
    .B(net27),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_4 c94 (.A(net985),
    .B(net820),
    .Y(net31));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net820),
    .B(net847),
    .Y(net32));
 sky130_fd_sc_hd__xnor2_4 c96 (.A(net27),
    .B(net25),
    .Y(net33));
 sky130_fd_sc_hd__xnor2_2 c97 (.A(net14),
    .B(net834),
    .Y(net34));
 sky130_fd_sc_hd__a41o_1 c98 (.A1(net28),
    .A2(net834),
    .A3(net869),
    .A4(net860),
    .B1(net32),
    .X(net35));
 sky130_fd_sc_hd__a21bo_2 c99 (.A1(net6),
    .A2(net28),
    .B1_N(net31),
    .X(net36));
 sky130_fd_sc_hd__a31o_1 merge763 (.A1(net406),
    .A2(net64),
    .A3(net404),
    .B1(clknet_1_0__leaf_net516),
    .X(net627));
 sky130_fd_sc_hd__a31o_1 merge764 (.A1(net51),
    .A2(net36),
    .A3(net50),
    .B1(net932),
    .X(net628));
 sky130_fd_sc_hd__a31o_1 merge765 (.A1(net822),
    .A2(net295),
    .A3(net296),
    .B1(net192),
    .X(net629));
 sky130_fd_sc_hd__a31o_1 merge766 (.A1(net106),
    .A2(net111),
    .A3(net113),
    .B1(net943),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 merge767 (.A0(net230),
    .A1(net133),
    .A2(net862),
    .A3(net254),
    .S0(net970),
    .S1(clknet_1_0__leaf_net919),
    .X(net631));
 sky130_fd_sc_hd__a31o_1 merge768 (.A1(net86),
    .A2(net100),
    .A3(net95),
    .B1(net91),
    .X(net632));
 sky130_fd_sc_hd__a31o_1 merge769 (.A1(net296),
    .A2(net200),
    .A3(net408),
    .B1(net402),
    .X(net633));
 sky130_fd_sc_hd__a31o_1 merge770 (.A1(net215),
    .A2(net949),
    .A3(net222),
    .B1(net308),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 merge771 (.A0(net152),
    .A1(net61),
    .A2(net925),
    .A3(net170),
    .S0(net928),
    .S1(net840),
    .X(net635));
 sky130_fd_sc_hd__a41o_1 merge772 (.A1(net219),
    .A2(net123),
    .A3(net128),
    .A4(net937),
    .B1(net91),
    .X(net636));
 sky130_fd_sc_hd__a31o_1 merge773 (.A1(net135),
    .A2(net155),
    .A3(clknet_1_0__leaf_net158),
    .B1(net159),
    .X(net637));
 sky130_fd_sc_hd__sdfrtp_1 merge774 (.CLK(clknet_4_4_0_clk),
    .D(net411),
    .RESET_B(clknet_1_1__leaf_net327),
    .SCD(net437),
    .SCE(net426),
    .Q(net638));
 sky130_fd_sc_hd__mux4_1 merge775 (.A0(net131),
    .A1(net117),
    .A2(net944),
    .A3(net863),
    .S0(net114),
    .S1(net135),
    .X(net639));
 sky130_fd_sc_hd__a41o_1 merge776 (.A1(net315),
    .A2(net235),
    .A3(net241),
    .A4(net319),
    .B1(net323),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net215),
    .A1(net206),
    .A2(net835),
    .A3(net222),
    .S0(net221),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net356),
    .A1(net403),
    .A2(net409),
    .A3(net338),
    .S0(net231),
    .S1(net449),
    .X(net642));
 sky130_fd_sc_hd__a41o_1 merge779 (.A1(net849),
    .A2(net263),
    .A3(net254),
    .A4(net271),
    .B1(net269),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(clknet_1_1__leaf_net327),
    .A1(net208),
    .A2(net201),
    .A3(net430),
    .S0(net426),
    .S1(net945),
    .X(net644));
 sky130_fd_sc_hd__a31o_1 merge781 (.A1(clknet_1_0__leaf_net516),
    .A2(net945),
    .A3(net408),
    .B1(net415),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_1 merge782 (.A(net700),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net1028),
    .A1(net119),
    .A2(net130),
    .A3(net141),
    .S0(net1029),
    .S1(net1000),
    .X(net647));
 sky130_fd_sc_hd__a41o_1 merge784 (.A1(net159),
    .A2(net152),
    .A3(net144),
    .A4(net82),
    .B1(net938),
    .X(net648));
 sky130_fd_sc_hd__mux4_1 merge785 (.A0(net54),
    .A1(net60),
    .A2(net856),
    .A3(net171),
    .S0(net960),
    .S1(net1015),
    .X(net649));
 sky130_fd_sc_hd__sdfbbn_1 merge786 (.CLK_N(clknet_4_1_0_clk),
    .D(net317),
    .RESET_B(net305),
    .SCD(net440),
    .SCE(net437),
    .SET_B(net434),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__mux4_1 merge787 (.A0(net46),
    .A1(net50),
    .A2(net56),
    .A3(net921),
    .S0(net60),
    .S1(net1014),
    .X(net652));
 sky130_fd_sc_hd__mux4_1 merge788 (.A0(net345),
    .A1(net338),
    .A2(net899),
    .A3(net296),
    .S0(net291),
    .S1(net818),
    .X(net653));
 sky130_fd_sc_hd__mux4_1 merge789 (.A0(net831),
    .A1(net937),
    .A2(net67),
    .A3(net305),
    .S0(net291),
    .S1(net321),
    .X(net654));
 sky130_fd_sc_hd__mux4_1 merge790 (.A0(net346),
    .A1(net358),
    .A2(clknet_1_0__leaf_net329),
    .A3(net899),
    .S0(net688),
    .S1(net763),
    .X(net655));
 sky130_fd_sc_hd__mux4_1 merge791 (.A0(net313),
    .A1(clknet_1_0__leaf_net327),
    .A2(net324),
    .A3(net409),
    .S0(net403),
    .S1(net405),
    .X(net656));
 sky130_fd_sc_hd__a31o_1 merge792 (.A1(net422),
    .A2(net415),
    .A3(net526),
    .B1(net1016),
    .X(net657));
 sky130_fd_sc_hd__a31o_1 merge793 (.A1(clknet_1_1__leaf_net516),
    .A2(net529),
    .A3(net64),
    .B1(net422),
    .X(net658));
 sky130_fd_sc_hd__a41o_1 merge794 (.A1(net426),
    .A2(net412),
    .A3(clknet_1_0__leaf_net327),
    .A4(net319),
    .B1(net667),
    .X(net659));
 sky130_fd_sc_hd__mux4_1 merge795 (.A0(net208),
    .A1(clknet_1_1__leaf_net327),
    .A2(net405),
    .A3(net532),
    .S0(net412),
    .S1(net535),
    .X(net660));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net415),
    .A1(net412),
    .A2(net187),
    .A3(net534),
    .S0(net522),
    .S1(net533),
    .X(net661));
 sky130_fd_sc_hd__a41o_1 merge797 (.A1(net418),
    .A2(net415),
    .A3(net294),
    .A4(net292),
    .B1(net200),
    .X(net662));
 sky130_fd_sc_hd__dfrbp_1 merge798 (.CLK(clknet_4_1_0_clk),
    .D(net629),
    .RESET_B(net310),
    .Q(net664),
    .Q_N(net663));
 sky130_fd_sc_hd__dfrbp_1 merge799 (.CLK(clknet_4_11_0_clk),
    .D(net384),
    .RESET_B(net388),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__dfrtn_1 merge800 (.CLK_N(clknet_4_0_0_clk),
    .D(net330),
    .RESET_B(net634),
    .Q(net667));
 sky130_fd_sc_hd__dfrtp_1 merge801 (.CLK(clknet_4_2_0_clk),
    .D(net630),
    .RESET_B(net647),
    .Q(net668));
 sky130_fd_sc_hd__dfrtp_1 merge802 (.CLK(clknet_4_2_0_clk),
    .D(net212),
    .Q(net641));
 sky130_fd_sc_hd__dfrtp_2 merge803 (.CLK(clknet_4_8_0_clk),
    .D(net156),
    .RESET_B(net637),
    .Q(net670));
 sky130_fd_sc_hd__dfsbp_1 merge804 (.CLK(clknet_4_11_0_clk),
    .SET_B(net289),
    .Q(net924),
    .Q_N(net290));
 sky130_fd_sc_hd__xnor2_1 merge805 (.A(net566),
    .B(net574),
    .Y(net672));
 sky130_fd_sc_hd__dfsbp_1 merge806 (.CLK(clknet_4_5_0_clk),
    .D(net551),
    .SET_B(net556),
    .Q(net674),
    .Q_N(net673));
 sky130_fd_sc_hd__dfstp_1 merge807 (.CLK(clknet_4_11_0_clk),
    .D(net286),
    .SET_B(net631),
    .Q(net675));
 sky130_fd_sc_hd__dfstp_1 merge808 (.CLK(clknet_4_4_0_clk),
    .D(net633),
    .SET_B(net661),
    .Q(net676));
 sky130_fd_sc_hd__dfstp_1 merge809 (.CLK(clknet_4_4_0_clk),
    .D(net443),
    .SET_B(net442),
    .Q(net677));
 sky130_fd_sc_hd__dlrbn_1 merge810 (.D(net628),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net649),
    .Q(net679),
    .Q_N(net678));
 sky130_fd_sc_hd__dlrbn_1 merge811 (.D(net250),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net257),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dlrbp_1 merge812 (.D(net527),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net627),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net178),
    .B(net180),
    .Y(net684));
 sky130_fd_sc_hd__dlrbp_1 merge814 (.D(net361),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net364),
    .Q(net686),
    .Q_N(net685));
 sky130_fd_sc_hd__dlrtn_1 merge815 (.D(net232),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net234),
    .Q(net687));
 sky130_fd_sc_hd__dlrtn_1 merge816 (.D(net339),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net342),
    .Q(net688));
 sky130_fd_sc_hd__dlrtn_1 merge817 (.D(net485),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net470),
    .Q(net689));
 sky130_fd_sc_hd__dlrtp_1 merge818 (.D(net499),
    .GATE(clknet_4_15_0_clk),
    .Q(net500));
 sky130_fd_sc_hd__xnor2_1 merge819 (.A(net136),
    .B(net145),
    .Y(net691));
 sky130_fd_sc_hd__dlrtp_1 merge820 (.D(net632),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net104),
    .Q(net692));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net626),
    .B(net612),
    .Y(net693));
 sky130_fd_sc_hd__dlrtp_1 merge822 (.D(net466),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net452),
    .Q(net694));
 sky130_fd_sc_hd__edfxbp_1 merge823 (.CLK(clknet_4_7_0_clk),
    .D(net589),
    .DE(net590),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__xnor2_1 merge824 (.A(net558),
    .B(net610),
    .Y(net697));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net576),
    .B(net508),
    .Y(net698));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net149),
    .B(net377),
    .Y(net699));
 sky130_fd_sc_hd__edfxtp_1 merge827 (.CLK(clknet_4_4_0_clk),
    .D(net662),
    .DE(net645),
    .Q(net700));
 sky130_fd_sc_hd__sdlclkp_1 merge828 (.CLK(clknet_4_9_0_clk),
    .GATE(net243),
    .SCE(net247),
    .GCLK(net701));
 sky130_fd_sc_hd__xnor2_1 merge829 (.A(net181),
    .B(net183),
    .Y(net702));
 sky130_fd_sc_hd__sdlclkp_2 merge830 (.CLK(clknet_4_10_0_clk),
    .GATE(net702),
    .SCE(net684),
    .GCLK(net891));
 sky130_fd_sc_hd__sdlclkp_4 merge831 (.CLK(clknet_4_6_0_clk),
    .GATE(net468),
    .SCE(net698),
    .GCLK(net703));
 sky130_fd_sc_hd__dfrbp_1 merge832 (.CLK(clknet_4_4_0_clk),
    .D(net656),
    .RESET_B(net660),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__dfrbp_1 merge833 (.CLK(clknet_4_1_0_clk),
    .D(net653),
    .RESET_B(net654),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dfrtn_1 merge834 (.CLK_N(clknet_4_8_0_clk),
    .D(net639),
    .RESET_B(net648),
    .Q(net708));
 sky130_fd_sc_hd__dfrtp_1 merge835 (.CLK(clknet_4_13_0_clk),
    .D(net597),
    .RESET_B(net625),
    .Q(net709));
 sky130_fd_sc_hd__dfrtp_1 merge836 (.CLK(clknet_4_15_0_clk),
    .D(net595),
    .RESET_B(net624),
    .Q(net710));
 sky130_fd_sc_hd__dfrtp_1 merge837 (.CLK(clknet_4_0_0_clk),
    .RESET_B(net218),
    .Q(net224));
 sky130_fd_sc_hd__dfsbp_1 merge838 (.CLK(clknet_4_7_0_clk),
    .D(net608),
    .SET_B(net599),
    .Q(net713),
    .Q_N(net712));
 sky130_fd_sc_hd__dfsbp_1 merge839 (.CLK(clknet_4_8_0_clk),
    .D(net691),
    .SET_B(net699),
    .Q(net715),
    .Q_N(net714));
 sky130_fd_sc_hd__xnor2_1 merge840 (.A(net400),
    .B(net399),
    .Y(net716));
 sky130_fd_sc_hd__dfstp_1 merge841 (.CLK(clknet_4_2_0_clk),
    .D(net118),
    .Q(net120));
 sky130_fd_sc_hd__dfstp_1 merge842 (.CLK(clknet_4_12_0_clk),
    .D(net370),
    .SET_B(net514),
    .Q(net718));
 sky130_fd_sc_hd__dfstp_1 merge843 (.CLK(clknet_4_5_0_clk),
    .D(net697),
    .SET_B(net658),
    .Q(net719));
 sky130_fd_sc_hd__dlrbn_1 merge844 (.D(net672),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net657),
    .Q(net721),
    .Q_N(net720));
 sky130_fd_sc_hd__dlrbn_1 merge845 (.D(net640),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net659),
    .Q(net723),
    .Q_N(net722));
 sky130_fd_sc_hd__dlrbp_1 merge846 (.D(net373),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net621),
    .Q(net725),
    .Q_N(net724));
 sky130_fd_sc_hd__dlrbp_1 merge847 (.D(net643),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net636),
    .Q(net727),
    .Q_N(net726));
 sky130_fd_sc_hd__dlrtn_1 merge848 (.D(net635),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net652),
    .Q(net728));
 sky130_fd_sc_hd__dlrtn_1 merge849 (.D(net454),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net492),
    .Q(net729));
 sky130_fd_sc_hd__xnor2_1 merge850 (.A(net395),
    .B(net716),
    .Y(net730));
 sky130_fd_sc_hd__xnor2_1 merge851 (.A(net392),
    .B(net509),
    .Y(net731));
 sky130_fd_sc_hd__dlrtn_2 merge852 (.D(net731),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net264),
    .Q(net898));
 sky130_fd_sc_hd__dlrtp_1 merge853 (.D(net613),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net614),
    .Q(net732));
 sky130_fd_sc_hd__dlrtp_1 merge854 (.D(net40),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net265),
    .Q(net932));
 sky130_fd_sc_hd__dlrtp_1 merge855 (.D(net693),
    .GATE(clknet_4_15_0_clk),
    .Q(net733));
 sky130_fd_sc_hd__edfxbp_1 merge856 (.CLK(clknet_4_14_0_clk),
    .D(net730),
    .DE(net362),
    .Q(net910),
    .Q_N(net734));
 sky130_fd_sc_hd__dfxbp_1 s857 (.CLK(clknet_4_10_0_clk),
    .D(net59),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__dfxbp_1 s858 (.CLK(clknet_4_10_0_clk),
    .D(net63),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dfxtp_2 s859 (.CLK(clknet_4_2_0_clk),
    .D(net126),
    .Q(net739));
 sky130_fd_sc_hd__dfxtp_1 s860 (.CLK(clknet_4_8_0_clk),
    .D(net142),
    .Q(net740));
 sky130_fd_sc_hd__dfxtp_2 s861 (.CLK(clknet_4_8_0_clk),
    .D(net143),
    .Q(net741));
 sky130_fd_sc_hd__dlclkp_1 s862 (.CLK(clknet_4_8_0_clk),
    .GATE(net150),
    .GCLK(net742));
 sky130_fd_sc_hd__dlclkp_2 s863 (.CLK(clknet_4_8_0_clk),
    .GATE(net157),
    .GCLK(net743));
 sky130_fd_sc_hd__dlclkp_4 s864 (.CLK(clknet_4_10_0_clk),
    .GATE(net163),
    .GCLK(net919));
 sky130_fd_sc_hd__dlxbn_2 s865 (.D(net164),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net745),
    .Q_N(net744));
 sky130_fd_sc_hd__dlxbn_1 s866 (.D(net166),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net927),
    .Q_N(net746));
 sky130_fd_sc_hd__dlxbp_1 s867 (.D(net169),
    .GATE(clknet_4_10_0_clk),
    .Q(net920),
    .Q_N(net747));
 sky130_fd_sc_hd__dlxtn_1 s868 (.D(net177),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net748));
 sky130_fd_sc_hd__dlxtn_1 s869 (.D(net182),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net903));
 sky130_fd_sc_hd__dlxtn_4 s870 (.D(net204),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net749));
 sky130_fd_sc_hd__dlxtp_1 s871 (.D(net210),
    .GATE(clknet_4_0_0_clk),
    .Q(net750));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s872 (.D(net225),
    .SLEEP_B(clknet_4_2_0_clk),
    .Q(net751));
 sky130_fd_sc_hd__dfxbp_1 s873 (.CLK(clknet_4_2_0_clk),
    .D(net238),
    .Q(net753),
    .Q_N(net752));
 sky130_fd_sc_hd__dfxbp_1 s874 (.CLK(clknet_4_9_0_clk),
    .D(net245),
    .Q(net755),
    .Q_N(net754));
 sky130_fd_sc_hd__dfxtp_1 s875 (.CLK(clknet_4_3_0_clk),
    .D(net246),
    .Q(net756));
 sky130_fd_sc_hd__dfxtp_1 s876 (.CLK(clknet_4_9_0_clk),
    .D(net267),
    .Q(net757));
 sky130_fd_sc_hd__dfxtp_1 s877 (.CLK(clknet_4_9_0_clk),
    .D(net279),
    .Q(net758));
 sky130_fd_sc_hd__dlclkp_1 s878 (.CLK(clknet_4_11_0_clk),
    .GATE(net288),
    .GCLK(net906));
 sky130_fd_sc_hd__dlclkp_2 s879 (.CLK(clknet_4_1_0_clk),
    .GATE(net311),
    .GCLK(net759));
 sky130_fd_sc_hd__dlclkp_4 s880 (.CLK(clknet_4_0_0_clk),
    .GATE(net325),
    .GCLK(net760));
 sky130_fd_sc_hd__dlxbn_1 s881 (.D(net332),
    .GATE_N(clknet_4_4_0_clk),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__dlxbn_1 s882 (.D(net341),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__dlxbp_1 s883 (.D(net351),
    .GATE(clknet_4_3_0_clk),
    .Q(net766),
    .Q_N(net765));
 sky130_fd_sc_hd__dlxtn_2 s884 (.D(net367),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net767));
 sky130_fd_sc_hd__dlxtn_1 s885 (.D(net369),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net768));
 sky130_fd_sc_hd__dlxtn_1 s886 (.D(net374),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net888));
 sky130_fd_sc_hd__dlxtp_1 s887 (.D(net376),
    .GATE(clknet_4_14_0_clk),
    .Q(net900));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s888 (.D(net380),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net769));
 sky130_fd_sc_hd__dfxbp_1 s889 (.CLK(clknet_4_11_0_clk),
    .D(net389),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__dfxbp_1 s890 (.CLK(clknet_4_11_0_clk),
    .D(net391),
    .Q(net773),
    .Q_N(net772));
 sky130_fd_sc_hd__dfxtp_1 s891 (.CLK(clknet_4_11_0_clk),
    .D(net396),
    .Q(net774));
 sky130_fd_sc_hd__dfxtp_2 s892 (.CLK(clknet_4_4_0_clk),
    .D(net423),
    .Q(net775));
 sky130_fd_sc_hd__dfxtp_2 s893 (.CLK(clknet_4_4_0_clk),
    .D(net433),
    .Q(net776));
 sky130_fd_sc_hd__dlclkp_1 s894 (.CLK(clknet_4_6_0_clk),
    .GATE(net459),
    .GCLK(net777));
 sky130_fd_sc_hd__dlclkp_2 s895 (.CLK(clknet_4_3_0_clk),
    .GATE(net460),
    .GCLK(net778));
 sky130_fd_sc_hd__dlclkp_4 s896 (.CLK(clknet_4_6_0_clk),
    .GATE(net463),
    .GCLK(net779));
 sky130_fd_sc_hd__dlxbn_1 s897 (.D(net464),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dlxbn_1 s898 (.D(net465),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net783),
    .Q_N(net782));
 sky130_fd_sc_hd__dlxbp_1 s899 (.D(net467),
    .GATE(clknet_4_6_0_clk),
    .Q(net785),
    .Q_N(net784));
 sky130_fd_sc_hd__dlxtn_1 s900 (.D(net469),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net786));
 sky130_fd_sc_hd__dlxtn_1 s901 (.D(net480),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net935));
 sky130_fd_sc_hd__dlxtn_1 s902 (.D(net483),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net787));
 sky130_fd_sc_hd__dlxtp_1 s903 (.D(net484),
    .GATE(clknet_4_12_0_clk),
    .Q(net788));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s904 (.D(net486),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net885));
 sky130_fd_sc_hd__dfxbp_1 s905 (.CLK(clknet_4_6_0_clk),
    .D(net487),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__dfxbp_1 s906 (.CLK(clknet_4_13_0_clk),
    .D(net488),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__dfxtp_1 s907 (.CLK(clknet_4_13_0_clk),
    .D(net490),
    .Q(net793));
 sky130_fd_sc_hd__dfxtp_1 s908 (.CLK(clknet_4_15_0_clk),
    .D(net494),
    .Q(net794));
 sky130_fd_sc_hd__dfxtp_1 s909 (.CLK(clknet_4_14_0_clk),
    .D(net504),
    .Q(net795));
 sky130_fd_sc_hd__dlclkp_1 s910 (.CLK(clknet_4_5_0_clk),
    .GATE(net560),
    .GCLK(net796));
 sky130_fd_sc_hd__dlclkp_2 s911 (.CLK(clknet_4_5_0_clk),
    .GATE(net575),
    .GCLK(net797));
 sky130_fd_sc_hd__dlclkp_4 s912 (.CLK(clknet_4_5_0_clk),
    .GATE(net577),
    .GCLK(net798));
 sky130_fd_sc_hd__dlxbn_1 s913 (.D(net579),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net800),
    .Q_N(net799));
 sky130_fd_sc_hd__dlxbn_1 s914 (.D(net583),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net802),
    .Q_N(net801));
 sky130_fd_sc_hd__dlxbp_1 s915 (.D(net584),
    .GATE(clknet_4_7_0_clk),
    .Q(net804),
    .Q_N(net803));
 sky130_fd_sc_hd__dlxtn_2 s916 (.D(net587),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net805));
 sky130_fd_sc_hd__dlxtn_1 s917 (.D(net588),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net806));
 sky130_fd_sc_hd__dlxtn_1 s918 (.D(net593),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net807));
 sky130_fd_sc_hd__dlxtp_1 s919 (.D(net609),
    .GATE(clknet_4_13_0_clk),
    .Q(net808));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s920 (.D(net615),
    .SLEEP_B(clknet_4_15_0_clk),
    .Q(net809));
 sky130_fd_sc_hd__dfxbp_1 s921 (.CLK(clknet_4_15_0_clk),
    .D(net616),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__dfxbp_1 s922 (.CLK(clknet_4_13_0_clk),
    .D(net619),
    .Q(net813),
    .Q_N(net812));
 sky130_fd_sc_hd__dfxtp_1 s923 (.CLK(clknet_4_3_0_clk),
    .D(net642),
    .Q(net814));
 sky130_fd_sc_hd__dfxtp_1 s924 (.CLK(clknet_4_4_0_clk),
    .D(net644),
    .Q(net815));
 sky130_fd_sc_hd__dfxtp_1 s925 (.CLK(clknet_4_12_0_clk),
    .D(net655),
    .Q(net816));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(in0),
    .X(net618));
 sky130_fd_sc_hd__buf_2 input2 (.A(in1),
    .X(net671));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net817));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net819));
 sky130_fd_sc_hd__buf_6 input6 (.A(in13),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(in16),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(in17),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(in18),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net826));
 sky130_fd_sc_hd__buf_6 input13 (.A(in2),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(in21),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in22),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net831));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in24),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in25),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net834));
 sky130_fd_sc_hd__buf_6 input21 (.A(in27),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in28),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net838));
 sky130_fd_sc_hd__buf_1 input25 (.A(in30),
    .X(net839));
 sky130_fd_sc_hd__buf_4 input26 (.A(in31),
    .X(net840));
 sky130_fd_sc_hd__buf_1 input27 (.A(in32),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input28 (.A(in33),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in34),
    .X(net843));
 sky130_fd_sc_hd__buf_1 input30 (.A(in35),
    .X(net844));
 sky130_fd_sc_hd__buf_8 input31 (.A(in36),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in37),
    .X(net846));
 sky130_fd_sc_hd__buf_4 input33 (.A(in38),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input34 (.A(in39),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(in4),
    .X(net849));
 sky130_fd_sc_hd__buf_1 input36 (.A(in40),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(in41),
    .X(net851));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input39 (.A(in43),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in44),
    .X(net854));
 sky130_fd_sc_hd__buf_2 input41 (.A(in45),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(in46),
    .X(net856));
 sky130_fd_sc_hd__buf_1 input43 (.A(in47),
    .X(net857));
 sky130_fd_sc_hd__dlymetal6s2s_1 input44 (.A(in48),
    .X(net858));
 sky130_fd_sc_hd__buf_1 input45 (.A(in49),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(in5),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(in50),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in51),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in52),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in53),
    .X(net864));
 sky130_fd_sc_hd__buf_4 input51 (.A(in54),
    .X(net865));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(in56),
    .X(net867));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net869));
 sky130_fd_sc_hd__buf_2 input56 (.A(in59),
    .X(net870));
 sky130_fd_sc_hd__buf_4 input57 (.A(in6),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(in60),
    .X(net872));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(in7),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in8),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_8 input62 (.A(in9),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net877),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net878),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output65 (.A(net879),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output66 (.A(net880),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output67 (.A(net881),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output68 (.A(net882),
    .X(out14));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net883),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output70 (.A(net884),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output71 (.A(net885),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output72 (.A(net886),
    .X(out18));
 sky130_fd_sc_hd__buf_2 output73 (.A(net887),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output74 (.A(net888),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(clknet_1_1__leaf_net889),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output76 (.A(net890),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(clknet_1_1__leaf_net891),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output78 (.A(net892),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output79 (.A(net893),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output80 (.A(net894),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output81 (.A(net895),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output82 (.A(net896),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output83 (.A(net897),
    .X(out29));
 sky130_fd_sc_hd__buf_2 output84 (.A(net898),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output85 (.A(net899),
    .X(out30));
 sky130_fd_sc_hd__buf_2 output86 (.A(net900),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output87 (.A(net901),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(clknet_1_0__leaf_net902),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output89 (.A(net903),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output90 (.A(net904),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output91 (.A(net905),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(clknet_1_1__leaf_net906),
    .X(out37));
 sky130_fd_sc_hd__buf_2 output93 (.A(net907),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output94 (.A(net908),
    .X(out39));
 sky130_fd_sc_hd__buf_2 output95 (.A(net909),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output96 (.A(net910),
    .X(out40));
 sky130_fd_sc_hd__buf_2 output97 (.A(net944),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output98 (.A(net912),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output99 (.A(net960),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output100 (.A(net914),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output101 (.A(net915),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output102 (.A(net916),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output103 (.A(net917),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output104 (.A(net918),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(clknet_1_1__leaf_net919),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output106 (.A(net920),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output107 (.A(net921),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output108 (.A(net922),
    .X(out51));
 sky130_fd_sc_hd__buf_2 output109 (.A(net923),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output110 (.A(net924),
    .X(out53));
 sky130_fd_sc_hd__buf_2 output111 (.A(net925),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output112 (.A(net926),
    .X(out55));
 sky130_fd_sc_hd__buf_2 output113 (.A(net927),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output114 (.A(net928),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output115 (.A(net929),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output116 (.A(net947),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output117 (.A(net931),
    .X(out60));
 sky130_fd_sc_hd__buf_2 output118 (.A(net932),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output119 (.A(net933),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output120 (.A(net934),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output121 (.A(net935),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net477),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net105),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net29),
    .X(net938));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(net366),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net335),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(net229),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net115),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout130 (.A(net973),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net304),
    .X(net945));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net201),
    .X(net946));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net930),
    .X(net947));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(net930),
    .X(net948));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net87),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net227),
    .X(net952));
 sky130_fd_sc_hd__buf_8 fanout139 (.A(net878),
    .X(net953));
 sky130_fd_sc_hd__buf_8 fanout140 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__buf_8 fanout142 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_12 fanout143 (.A(net13),
    .X(net957));
 sky130_fd_sc_hd__buf_4 max_cap144 (.A(net76),
    .X(net958));
 sky130_fd_sc_hd__buf_4 max_cap145 (.A(net887),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net913),
    .X(net960));
 sky130_fd_sc_hd__buf_4 max_cap147 (.A(net69),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net769),
    .X(net962));
 sky130_fd_sc_hd__buf_2 max_cap149 (.A(net751),
    .X(net963));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net741),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net552),
    .X(net965));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(net553),
    .X(net966));
 sky130_fd_sc_hd__buf_4 max_cap153 (.A(net74),
    .X(net967));
 sky130_fd_sc_hd__buf_12 fanout154 (.A(net827),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net798 (.A(net798),
    .X(clknet_0_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_0__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net798 (.A(clknet_0_net798),
    .X(clknet_1_1__leaf_net798));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net797 (.A(net797),
    .X(clknet_0_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_0__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net797 (.A(clknet_0_net797),
    .X(clknet_1_1__leaf_net797));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net796 (.A(net796),
    .X(clknet_0_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_0__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net796 (.A(clknet_0_net796),
    .X(clknet_1_1__leaf_net796));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net591 (.A(net591),
    .X(clknet_0_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_0__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net591 (.A(clknet_0_net591),
    .X(clknet_1_1__leaf_net591));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net565 (.A(net565),
    .X(clknet_0_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_0__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net565 (.A(clknet_0_net565),
    .X(clknet_1_1__leaf_net565));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net779 (.A(net779),
    .X(clknet_0_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_0__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net779 (.A(clknet_0_net779),
    .X(clknet_1_1__leaf_net779));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net778 (.A(net778),
    .X(clknet_0_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net778 (.A(clknet_0_net778),
    .X(clknet_1_0__leaf_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net778 (.A(clknet_0_net778),
    .X(clknet_1_1__leaf_net778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net777 (.A(net777),
    .X(clknet_0_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_0__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net777 (.A(clknet_0_net777),
    .X(clknet_1_1__leaf_net777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net760 (.A(net760),
    .X(clknet_0_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net760 (.A(clknet_0_net760),
    .X(clknet_1_1__leaf_net760));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net479 (.A(net479),
    .X(clknet_0_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_0__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net479 (.A(clknet_0_net479),
    .X(clknet_1_1__leaf_net479));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net457 (.A(net457),
    .X(clknet_0_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_0__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net457 (.A(clknet_0_net457),
    .X(clknet_1_1__leaf_net457));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net458 (.A(net458),
    .X(clknet_0_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_0__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net458 (.A(clknet_0_net458),
    .X(clknet_1_1__leaf_net458));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net435 (.A(net435),
    .X(clknet_0_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_0__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net435 (.A(clknet_0_net435),
    .X(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net546 (.A(net546),
    .X(clknet_0_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_0__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net546 (.A(clknet_0_net546),
    .X(clknet_1_1__leaf_net546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net538 (.A(net538),
    .X(clknet_0_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_0__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net538 (.A(clknet_0_net538),
    .X(clknet_1_1__leaf_net538));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net703 (.A(net703),
    .X(clknet_0_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net471 (.A(net471),
    .X(clknet_0_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_0__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net471 (.A(clknet_0_net471),
    .X(clknet_1_1__leaf_net471));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net542 (.A(net542),
    .X(clknet_0_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_0__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_1__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net557 (.A(net557),
    .X(clknet_0_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_0__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net557 (.A(clknet_0_net557),
    .X(clknet_1_1__leaf_net557));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net559 (.A(net559),
    .X(clknet_0_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_0__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net559 (.A(clknet_0_net559),
    .X(clknet_1_1__leaf_net559));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net554 (.A(net554),
    .X(clknet_0_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_0__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net554 (.A(clknet_0_net554),
    .X(clknet_1_1__leaf_net554));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net889 (.A(net889),
    .X(clknet_0_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_0__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net889 (.A(clknet_0_net889),
    .X(clknet_1_1__leaf_net889));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net378 (.A(net378),
    .X(clknet_0_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_0__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net378 (.A(clknet_0_net378),
    .X(clknet_1_1__leaf_net378));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net906 (.A(net906),
    .X(clknet_0_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_0__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net906 (.A(clknet_0_net906),
    .X(clknet_1_1__leaf_net906));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net919 (.A(net919),
    .X(clknet_0_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_0__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net919 (.A(clknet_0_net919),
    .X(clknet_1_1__leaf_net919));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net891 (.A(net891),
    .X(clknet_0_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_0__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net891 (.A(clknet_0_net891),
    .X(clknet_1_1__leaf_net891));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net743 (.A(net743),
    .X(clknet_0_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_0__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net743 (.A(clknet_0_net743),
    .X(clknet_1_1__leaf_net743));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net162 (.A(net162),
    .X(clknet_0_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_0__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net162 (.A(clknet_0_net162),
    .X(clknet_1_1__leaf_net162));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net742 (.A(net742),
    .X(clknet_0_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_0__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net742 (.A(clknet_0_net742),
    .X(clknet_1_1__leaf_net742));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net256 (.A(net256),
    .X(clknet_0_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_0__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net256 (.A(clknet_0_net256),
    .X(clknet_1_1__leaf_net256));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net283 (.A(net283),
    .X(clknet_0_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_0__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net283 (.A(clknet_0_net283),
    .X(clknet_1_1__leaf_net283));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net262 (.A(net262),
    .X(clknet_0_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_0__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net262 (.A(clknet_0_net262),
    .X(clknet_1_1__leaf_net262));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net251 (.A(net251),
    .X(clknet_0_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_0__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net251 (.A(clknet_0_net251),
    .X(clknet_1_1__leaf_net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net701 (.A(net701),
    .X(clknet_0_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net258 (.A(net258),
    .X(clknet_0_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_0__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_1__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net244 (.A(net244),
    .X(clknet_0_net244));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net244 (.A(clknet_0_net244),
    .X(clknet_1_0__leaf_net244));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net244 (.A(clknet_0_net244),
    .X(clknet_1_1__leaf_net244));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net21),
    .A1(net20),
    .A2(net982),
    .A3(net856),
    .S0(net6),
    .S1(net995),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net23),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net971),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net911),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net911),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net24),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net975),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net994),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net22),
    .X(net978));
 sky130_fd_sc_hd__buf_6 rebuffer11 (.A(net1),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net20),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net980),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net14),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net14),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_4 clone16 (.A(net827),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net12),
    .X(net985));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer18 (.A(net985),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net986),
    .X(net987));
 sky130_fd_sc_hd__buf_8 rebuffer20 (.A(net956),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net988),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(net989),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net988),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net991),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net1033),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_1 clone27 (.A(net955),
    .X(net995));
 sky130_fd_sc_hd__buf_6 rebuffer28 (.A(net1),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net955),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net567),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net811),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net740),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net714),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net601),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net568),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net677),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net345),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net707),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net300),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net696),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net755),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net776),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net382),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net749),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net805),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net932),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net747),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net524),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net708),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net667),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net774),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net525),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net386),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net792),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net885),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net767),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net450),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net788),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net724),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net121),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net739),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net812),
    .X(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_DE (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCD (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SCE (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_SCD (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A3 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A4 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_Q (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A4 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_SET_B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_SCD (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A4 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_Y (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_SCE (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A4 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_Q_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_SET_B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_SCD (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_Q (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_Y (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_B1_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SET_B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_D (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SCD (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1_N (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_SCE (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1_N (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_Y (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_Y (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A4 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_B1_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_Y (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCD (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SCE (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_D (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1_N (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_X (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A3 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_X (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_X (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_D (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_D (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_B1_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B1_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B1_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_B1_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_Y (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A4 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A3 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Y (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_Y (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A4 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_Y (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_S1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_Q (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_SET_B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_RESET_B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_DE (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_B1_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B1_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SCD (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_SCD (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_X (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_X (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_A2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_S1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A3 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SET_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_B (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_Y (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_S0 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_SCE (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_SCE (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_Y (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_D (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_X (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_RESET_B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCE (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_D (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_Q_N (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_Q (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_RESET_B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_S1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_Q_N (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_SCE (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_X (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_RESET_B (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A4 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_Q_N (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_X (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_SCD (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_D (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_B1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SCD (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S0 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_X (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A0 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_SCE (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A3 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_B1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_X (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_RESET_B (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A4 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_B (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_X (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_RESET_B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A4 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_RESET_B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_X (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_Q_N (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_RESET_B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_Q (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_SET_B (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_SCD (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_SCD (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_X (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A3 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_Q_N (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A3 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_Y (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_Q (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B1_N (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_Q (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A4 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A4 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_B1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_Q (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_Q (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_Q (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S1 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_RESET_B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q_N (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_B1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A4 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_Q (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_S1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_s870_Q (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_B (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_B1_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_Y (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_Q (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A4 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S1 (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1_N (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_Q (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A4 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1_N (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net759_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_GCLK (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_Y (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_Q_N (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SCE (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_B1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_Q (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_SCD (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_B1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_s884_Q (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_B1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCE (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_Q (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_B1_N (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_Q (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_SCE (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A4 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_B1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_Q (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_B1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_Q (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A4 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A4 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B1_N (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_Y (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_SCE (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_RESET_B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1_N (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A4 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_SCD (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1_N (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_B1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_S0 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_D (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1_N (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A3 (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A4 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_SCD (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1_N (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_B1_N (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A2 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A4 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_B1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_SCE (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1_N (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_B1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A4 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SCE (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A2 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A3 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A4 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SCD (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B1_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A3 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_S0 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_D (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_Y (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_S0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_Y (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_Q (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_Q (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_Q (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap145_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SCD (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_Y (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_Q (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_SET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_Y (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_Q (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A3 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A2 (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_Q (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_B1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_SET_B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_DE (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A4 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCD (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A3 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_S1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_SET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_Q (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_SCE (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_Q (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_Y (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_Q (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_RESET_B (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1_N (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_SCE (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_Q (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_Q (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_X (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A4 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_RESET_B (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_DE (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A4 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S0 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_D (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_B1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A0 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SET_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_SCE (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_SET_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_S0 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1_N (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_SET_B (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SET_B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A4 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_SET_B (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_D (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A4 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_B1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B1_N (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1_N (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_B1_N (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A4 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCE (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B1_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B1_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B1_N (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S0 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A4 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_RESET_B (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B1 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1_N (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1_N (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A4 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_RESET_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_B (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_B1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_D (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_SCD (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_X (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_B1 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap145_X (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A4 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_S1 (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_S0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_RESET_B (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap147_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_S1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A4 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_B1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A4 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A4 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A4 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_SCE (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_S0 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1_N (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_S1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_SCD (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A4 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_SCE (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_SCE (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A4 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_SCD (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_B1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s879_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s872_SLEEP_B (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s873_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s893_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s894_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s914_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_GATE (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_GATE_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s864_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s865_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s866_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s868_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s889_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s890_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s891_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_SLEEP_B (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_S1 (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B1 (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B1_N (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_SCE (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net760_X (.DIODE(clknet_1_0__leaf_net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net435_X (.DIODE(clknet_1_1__leaf_net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A2 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S1 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_RESET_B (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net363_X (.DIODE(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_SCD (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net363_X (.DIODE(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B1_N (.DIODE(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_B (.DIODE(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B1 (.DIODE(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net759_X (.DIODE(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_SET_B (.DIODE(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net759_X (.DIODE(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_S0 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A4 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_B1_N (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_S0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_SCE (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_RESET_B (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone25_X (.DIODE(net993));
 sky130_fd_sc_hd__clkbuf_1 clone1 (.A(net13),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_1 clone3 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net366),
    .X(net1033));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
