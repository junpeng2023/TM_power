module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net635;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net737;
 wire clknet_1_0__leaf_net737;
 wire clknet_1_1__leaf_net737;
 wire clknet_0_net592;
 wire clknet_1_0__leaf_net592;
 wire clknet_1_1__leaf_net592;
 wire clknet_0_net594;
 wire clknet_1_0__leaf_net594;
 wire clknet_1_1__leaf_net594;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net736;
 wire clknet_1_0__leaf_net736;
 wire clknet_1_1__leaf_net736;
 wire clknet_0_net719;
 wire clknet_1_0__leaf_net719;
 wire clknet_1_1__leaf_net719;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net480;
 wire clknet_1_0__leaf_net480;
 wire clknet_1_1__leaf_net480;
 wire clknet_0_net478;
 wire clknet_1_0__leaf_net478;
 wire clknet_1_1__leaf_net478;
 wire clknet_0_net701;
 wire clknet_1_0__leaf_net701;
 wire clknet_1_1__leaf_net701;
 wire clknet_0_net683;
 wire clknet_1_0__leaf_net683;
 wire clknet_1_1__leaf_net683;
 wire clknet_0_net462;
 wire clknet_1_0__leaf_net462;
 wire clknet_1_1__leaf_net462;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net682;
 wire clknet_1_0__leaf_net682;
 wire clknet_1_1__leaf_net682;
 wire clknet_0_net485;
 wire clknet_1_0__leaf_net485;
 wire clknet_1_1__leaf_net485;
 wire clknet_0_net681;
 wire clknet_1_0__leaf_net681;
 wire clknet_1_1__leaf_net681;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;

 sky130_fd_sc_hd__xnor2_2 c100 (.A(net817),
    .B(net829),
    .Y(net31));
 sky130_fd_sc_hd__a21bo_4 c101 (.A1(net23),
    .A2(net30),
    .B1_N(net29),
    .X(net32));
 sky130_fd_sc_hd__xnor2_2 c102 (.A(net32),
    .B(net28),
    .Y(net33));
 sky130_fd_sc_hd__a21bo_2 c103 (.A1(net25),
    .A2(net14),
    .B1_N(net919),
    .X(net34));
 sky130_fd_sc_hd__xnor2_1 c104 (.A(net34),
    .B(net33),
    .Y(net35));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net773),
    .A2(net817),
    .B1_N(net32),
    .X(net36));
 sky130_fd_sc_hd__a31o_1 c106 (.A1(net35),
    .A2(net29),
    .A3(net811),
    .B1(net32),
    .X(net37));
 sky130_fd_sc_hd__xnor2_1 c107 (.A(net30),
    .B(net34),
    .Y(net38));
 sky130_fd_sc_hd__a21bo_1 c108 (.A1(net37),
    .A2(net35),
    .B1_N(net783),
    .X(net39));
 sky130_fd_sc_hd__dfbbn_1 c109 (.CLK_N(clknet_4_4_0_clk),
    .D(net38),
    .RESET_B(net39),
    .SET_B(net26),
    .Q(net41),
    .Q_N(net40));
 sky130_fd_sc_hd__xnor2_4 c110 (.A(net22),
    .B(net791),
    .Y(net841));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net5),
    .B(net919),
    .Y(net850));
 sky130_fd_sc_hd__a21bo_1 c112 (.A1(net776),
    .A2(net12),
    .B1_N(net779),
    .X(net42));
 sky130_fd_sc_hd__a21bo_4 c113 (.A1(net827),
    .A2(net29),
    .B1_N(net922),
    .X(net43));
 sky130_fd_sc_hd__xnor2_1 c114 (.A(net43),
    .B(net25),
    .Y(net44));
 sky130_fd_sc_hd__xnor2_1 c115 (.A(net33),
    .B(net841),
    .Y(net45));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net28),
    .B(net42),
    .Y(net46));
 sky130_fd_sc_hd__xnor2_1 c117 (.A(net12),
    .B(net22),
    .Y(net47));
 sky130_fd_sc_hd__xnor2_1 c118 (.A(net47),
    .B(net780),
    .Y(net48));
 sky130_fd_sc_hd__xnor2_1 c119 (.A(net43),
    .B(net791),
    .Y(net49));
 sky130_fd_sc_hd__xnor2_4 c120 (.A(net29),
    .B(net843),
    .Y(net50));
 sky130_fd_sc_hd__xnor2_1 c121 (.A(net48),
    .B(net50),
    .Y(net51));
 sky130_fd_sc_hd__a21bo_2 c122 (.A1(net36),
    .A2(net43),
    .B1_N(net47),
    .X(net52));
 sky130_fd_sc_hd__xnor2_4 c123 (.A(net52),
    .B(net43),
    .Y(net863));
 sky130_fd_sc_hd__a21bo_1 c124 (.A1(net51),
    .A2(net48),
    .B1_N(net863),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 c125 (.A(net671),
    .X(net54));
 sky130_fd_sc_hd__a41o_1 c126 (.A1(net39),
    .A2(net635),
    .A3(net50),
    .A4(net818),
    .B1(net863),
    .X(net55));
 sky130_fd_sc_hd__a31o_1 c127 (.A1(net54),
    .A2(net25),
    .A3(net856),
    .B1(net43),
    .X(net56));
 sky130_fd_sc_hd__a41o_1 c128 (.A1(net14),
    .A2(net3),
    .A3(net43),
    .A4(net46),
    .B1(net863),
    .X(net57));
 sky130_fd_sc_hd__sdfbbn_1 c129 (.CLK_N(clknet_4_5_0_clk),
    .D(net53),
    .RESET_B(net43),
    .SCD(net866),
    .SCE(net841),
    .SET_B(net863),
    .Q(net870),
    .Q_N(net58));
 sky130_fd_sc_hd__sdfbbn_1 c130 (.CLK_N(clknet_4_5_0_clk),
    .D(net776),
    .RESET_B(net57),
    .SCD(net56),
    .SCE(net863),
    .SET_B(net50),
    .Q(net874),
    .Q_N(net59));
 sky130_fd_sc_hd__a41o_1 c131 (.A1(net52),
    .A2(net863),
    .A3(net59),
    .A4(net841),
    .B1(net671),
    .X(net60));
 sky130_fd_sc_hd__xnor2_4 c132 (.A(net790),
    .B(net770),
    .Y(net61));
 sky130_fd_sc_hd__xnor2_4 c133 (.A(net781),
    .B(net812),
    .Y(net62));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net827),
    .B(net769),
    .Y(net63));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net778),
    .B(net772),
    .Y(net64));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net918),
    .B(net768),
    .Y(net65));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net914),
    .B(net62),
    .Y(net66));
 sky130_fd_sc_hd__xnor2_4 c138 (.A(net775),
    .B(net823),
    .Y(net67));
 sky130_fd_sc_hd__xnor2_4 c139 (.A(net915),
    .B(net780),
    .Y(net68));
 sky130_fd_sc_hd__a21bo_4 c140 (.A1(net775),
    .A2(net67),
    .B1_N(net778),
    .X(net69));
 sky130_fd_sc_hd__xnor2_4 c141 (.A(net772),
    .B(net812),
    .Y(net70));
 sky130_fd_sc_hd__a21bo_4 c142 (.A1(net827),
    .A2(net774),
    .B1_N(net773),
    .X(net71));
 sky130_fd_sc_hd__xnor2_4 c143 (.A(net71),
    .B(net64),
    .Y(net72));
 sky130_fd_sc_hd__xnor2_4 c144 (.A(net917),
    .B(net937),
    .Y(net73));
 sky130_fd_sc_hd__xnor2_4 c145 (.A(net774),
    .B(net68),
    .Y(net74));
 sky130_fd_sc_hd__xnor2_4 c146 (.A(net70),
    .B(net812),
    .Y(net75));
 sky130_fd_sc_hd__mux4_2 c147 (.A0(net75),
    .A1(net72),
    .A2(net823),
    .A3(net917),
    .S0(net812),
    .S1(net915),
    .X(net76));
 sky130_fd_sc_hd__xnor2_4 c148 (.A(net69),
    .B(net778),
    .Y(net77));
 sky130_fd_sc_hd__xnor2_4 c149 (.A(net957),
    .B(net812),
    .Y(net78));
 sky130_fd_sc_hd__xnor2_2 c150 (.A(net790),
    .B(net916),
    .Y(net79));
 sky130_fd_sc_hd__a21bo_4 c151 (.A1(net907),
    .A2(net909),
    .B1_N(net66),
    .X(net80));
 sky130_fd_sc_hd__a21bo_4 c152 (.A1(net909),
    .A2(net77),
    .B1_N(net635),
    .X(net81));
 sky130_fd_sc_hd__xnor2_4 c153 (.A(net81),
    .B(net912),
    .Y(net832));
 sky130_fd_sc_hd__xnor2_4 c154 (.A(net909),
    .B(net69),
    .Y(net82));
 sky130_fd_sc_hd__xnor2_4 c155 (.A(net901),
    .B(net914),
    .Y(net83));
 sky130_fd_sc_hd__xnor2_4 c156 (.A(net801),
    .B(net83),
    .Y(net84));
 sky130_fd_sc_hd__a41o_4 c157 (.A1(net74),
    .A2(net804),
    .A3(net66),
    .A4(net795),
    .B1(net920),
    .X(net85));
 sky130_fd_sc_hd__xnor2_4 c158 (.A(net783),
    .B(net786),
    .Y(net86));
 sky130_fd_sc_hd__xnor2_4 c159 (.A(net920),
    .B(net85),
    .Y(net87));
 sky130_fd_sc_hd__xnor2_4 c160 (.A(net83),
    .B(net777),
    .Y(net88));
 sky130_fd_sc_hd__a31o_4 c161 (.A1(net86),
    .A2(net805),
    .A3(net87),
    .B1(net921),
    .X(net89));
 sky130_fd_sc_hd__a21bo_2 c162 (.A1(net778),
    .A2(net924),
    .B1_N(net901),
    .X(net90));
 sky130_fd_sc_hd__a21bo_2 c163 (.A1(net799),
    .A2(net74),
    .B1_N(net920),
    .X(net91));
 sky130_fd_sc_hd__a41o_4 c164 (.A1(net997),
    .A2(net828),
    .A3(net924),
    .A4(net771),
    .B1(net782),
    .X(net92));
 sky130_fd_sc_hd__xnor2_4 c165 (.A(net1029),
    .B(net89),
    .Y(net93));
 sky130_fd_sc_hd__a31o_2 c166 (.A1(net66),
    .A2(net92),
    .A3(net908),
    .B1(net920),
    .X(net94));
 sky130_fd_sc_hd__xnor2_4 c167 (.A(net94),
    .B(net92),
    .Y(net95));
 sky130_fd_sc_hd__a41o_2 c168 (.A1(net90),
    .A2(net70),
    .A3(net924),
    .A4(net95),
    .B1(net785),
    .X(net96));
 sky130_fd_sc_hd__xnor2_4 c169 (.A(net87),
    .B(net93),
    .Y(net97));
 sky130_fd_sc_hd__a41o_2 c170 (.A1(net95),
    .A2(net68),
    .A3(net86),
    .A4(net85),
    .B1(net72),
    .X(net98));
 sky130_fd_sc_hd__a31o_2 c171 (.A1(net88),
    .A2(net85),
    .A3(net73),
    .B1(net920),
    .X(net99));
 sky130_fd_sc_hd__a41o_4 c172 (.A1(net97),
    .A2(net788),
    .A3(net64),
    .A4(net82),
    .B1(net798),
    .X(net100));
 sky130_fd_sc_hd__a31o_1 c173 (.A1(net889),
    .A2(net92),
    .A3(net786),
    .B1(net84),
    .X(net101));
 sky130_fd_sc_hd__xnor2_2 c174 (.A(net98),
    .B(net827),
    .Y(net102));
 sky130_fd_sc_hd__a41o_2 c175 (.A1(net99),
    .A2(net101),
    .A3(net98),
    .A4(net891),
    .B1(net798),
    .X(net103));
 sky130_fd_sc_hd__a21bo_2 c176 (.A1(net823),
    .A2(net99),
    .B1_N(net920),
    .X(net104));
 sky130_fd_sc_hd__a21bo_4 c177 (.A1(net104),
    .A2(net98),
    .B1_N(net924),
    .X(net105));
 sky130_fd_sc_hd__a21bo_2 c178 (.A1(net774),
    .A2(net778),
    .B1_N(net104),
    .X(net106));
 sky130_fd_sc_hd__xnor2_4 c179 (.A(net820),
    .B(net105),
    .Y(net107));
 sky130_fd_sc_hd__a21bo_2 c180 (.A1(net73),
    .A2(net95),
    .B1_N(net104),
    .X(net108));
 sky130_fd_sc_hd__xnor2_2 c181 (.A(net75),
    .B(net804),
    .Y(net109));
 sky130_fd_sc_hd__a21bo_1 c182 (.A1(net101),
    .A2(net822),
    .B1_N(net109),
    .X(net110));
 sky130_fd_sc_hd__a21bo_4 c183 (.A1(net78),
    .A2(net803),
    .B1_N(net780),
    .X(net111));
 sky130_fd_sc_hd__a31o_4 c184 (.A1(net107),
    .A2(net822),
    .A3(net821),
    .B1(net997),
    .X(net112));
 sky130_fd_sc_hd__a31o_2 c185 (.A1(net814),
    .A2(net73),
    .A3(net890),
    .B1(net924),
    .X(net113));
 sky130_fd_sc_hd__xnor2_4 c186 (.A(net108),
    .B(net111),
    .Y(net114));
 sky130_fd_sc_hd__a21bo_2 c187 (.A1(net114),
    .A2(net101),
    .B1_N(net112),
    .X(net115));
 sky130_fd_sc_hd__a31o_4 c188 (.A1(net0),
    .A2(net111),
    .A3(net86),
    .B1(net110),
    .X(net116));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net814),
    .A1(net110),
    .A2(net810),
    .A3(net808),
    .S0(net890),
    .S1(net920),
    .X(net867));
 sky130_fd_sc_hd__a31o_1 c190 (.A1(net115),
    .A2(net814),
    .A3(net114),
    .B1(net803),
    .X(net117));
 sky130_fd_sc_hd__a31o_4 c191 (.A1(net825),
    .A2(net116),
    .A3(net819),
    .B1(net887),
    .X(net118));
 sky130_fd_sc_hd__mux4_2 c192 (.A0(net117),
    .A1(net108),
    .A2(net118),
    .A3(net112),
    .S0(net917),
    .S1(net867),
    .X(net119));
 sky130_fd_sc_hd__a21bo_2 c193 (.A1(net1011),
    .A2(net867),
    .B1_N(net790),
    .X(net120));
 sky130_fd_sc_hd__a21bo_1 c194 (.A1(net104),
    .A2(net120),
    .B1_N(net1014),
    .X(net121));
 sky130_fd_sc_hd__a31o_1 c195 (.A1(net119),
    .A2(net120),
    .A3(net99),
    .B1(net114),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net890),
    .A1(net997),
    .A2(net104),
    .A3(net121),
    .S0(net795),
    .S1(net907),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net121),
    .A1(net809),
    .A2(net109),
    .A3(net112),
    .S0(net120),
    .X(net124));
 sky130_fd_sc_hd__a21bo_1 c198 (.A1(net94),
    .A2(net786),
    .B1_N(net9),
    .X(net125));
 sky130_fd_sc_hd__xnor2_2 c199 (.A(net803),
    .B(net117),
    .Y(net126));
 sky130_fd_sc_hd__a21bo_1 c200 (.A1(net789),
    .A2(net8),
    .B1_N(net19),
    .X(net127));
 sky130_fd_sc_hd__a41o_1 c201 (.A1(net791),
    .A2(net8),
    .A3(net104),
    .A4(net111),
    .B1(net920),
    .X(net128));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net17),
    .A2(net931),
    .B1_N(net891),
    .X(net129));
 sky130_fd_sc_hd__a21bo_1 c203 (.A1(net786),
    .A2(net775),
    .B1_N(net3),
    .X(net130));
 sky130_fd_sc_hd__a21bo_1 c204 (.A1(net924),
    .A2(net808),
    .B1_N(net922),
    .X(net131));
 sky130_fd_sc_hd__a21bo_1 c205 (.A1(net117),
    .A2(net13),
    .B1_N(net892),
    .X(net132));
 sky130_fd_sc_hd__a31o_2 c206 (.A1(net98),
    .A2(net125),
    .A3(net128),
    .B1(net921),
    .X(net133));
 sky130_fd_sc_hd__a21bo_1 c207 (.A1(net108),
    .A2(net128),
    .B1_N(net6),
    .X(net134));
 sky130_fd_sc_hd__xnor2_4 c208 (.A(net10),
    .B(net889),
    .Y(net135));
 sky130_fd_sc_hd__a21bo_1 c209 (.A1(net2),
    .A2(net133),
    .B1_N(net132),
    .X(net136));
 sky130_fd_sc_hd__a31o_1 c210 (.A1(net128),
    .A2(net789),
    .A3(net867),
    .B1(net62),
    .X(net137));
 sky130_fd_sc_hd__a21bo_1 c211 (.A1(net132),
    .A2(net773),
    .B1_N(net133),
    .X(net138));
 sky130_fd_sc_hd__a31o_1 c212 (.A1(net86),
    .A2(net138),
    .A3(net135),
    .B1(net137),
    .X(net139));
 sky130_fd_sc_hd__a31o_1 c213 (.A1(net8),
    .A2(net113),
    .A3(net112),
    .B1(net907),
    .X(net140));
 sky130_fd_sc_hd__a21bo_1 c214 (.A1(net133),
    .A2(net125),
    .B1_N(net111),
    .X(net141));
 sky130_fd_sc_hd__a31o_2 c215 (.A1(net141),
    .A2(net804),
    .A3(net113),
    .B1(net140),
    .X(net142));
 sky130_fd_sc_hd__a31o_1 c216 (.A1(net13),
    .A2(net10),
    .A3(net1009),
    .B1(net133),
    .X(net143));
 sky130_fd_sc_hd__buf_1 c217 (.A(net671),
    .X(net859));
 sky130_fd_sc_hd__a31o_2 c218 (.A1(net140),
    .A2(net94),
    .A3(net141),
    .B1(net138),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net127),
    .A1(net3),
    .A2(net129),
    .A3(net136),
    .S0(net139),
    .S1(net907),
    .X(net145));
 sky130_fd_sc_hd__a21bo_1 c220 (.A1(net3),
    .A2(net119),
    .B1_N(net675),
    .X(net146));
 sky130_fd_sc_hd__xnor2_1 c221 (.A(net99),
    .B(net901),
    .Y(net147));
 sky130_fd_sc_hd__clkbuf_1 c222 (.A(net659),
    .X(net148));
 sky130_fd_sc_hd__a21bo_1 c223 (.A1(net774),
    .A2(net27),
    .B1_N(net9),
    .X(net149));
 sky130_fd_sc_hd__a21bo_1 c224 (.A1(net119),
    .A2(net818),
    .B1_N(net134),
    .X(net150));
 sky130_fd_sc_hd__buf_1 c225 (.A(net659),
    .X(net151));
 sky130_fd_sc_hd__a21bo_1 c226 (.A1(net828),
    .A2(net866),
    .B1_N(net892),
    .X(net152));
 sky130_fd_sc_hd__a31o_1 c227 (.A1(net774),
    .A2(net115),
    .A3(net791),
    .B1(net41),
    .X(net153));
 sky130_fd_sc_hd__a21bo_1 c228 (.A1(net127),
    .A2(net785),
    .B1_N(net151),
    .X(net154));
 sky130_fd_sc_hd__xnor2_1 c229 (.A(net778),
    .B(net143),
    .Y(net155));
 sky130_fd_sc_hd__xnor2_2 c230 (.A(net95),
    .B(net2),
    .Y(net156));
 sky130_fd_sc_hd__a21bo_1 c231 (.A1(net151),
    .A2(net136),
    .B1_N(net799),
    .X(net157));
 sky130_fd_sc_hd__xnor2_2 c232 (.A(net153),
    .B(net0),
    .Y(net158));
 sky130_fd_sc_hd__a31o_1 c233 (.A1(net785),
    .A2(net31),
    .A3(net152),
    .B1(net158),
    .X(net159));
 sky130_fd_sc_hd__a21bo_1 c234 (.A1(net41),
    .A2(net801),
    .B1_N(net24),
    .X(net160));
 sky130_fd_sc_hd__xnor2_1 c235 (.A(net133),
    .B(net36),
    .Y(net161));
 sky130_fd_sc_hd__a31o_1 c236 (.A1(net152),
    .A2(net896),
    .A3(net772),
    .B1(net867),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c237 (.A1(net154),
    .A2(net158),
    .B1_N(net159),
    .X(net163));
 sky130_fd_sc_hd__a41o_1 c238 (.A1(net27),
    .A2(net160),
    .A3(net32),
    .A4(net892),
    .B1(net24),
    .X(net835));
 sky130_fd_sc_hd__a21bo_1 c239 (.A1(net138),
    .A2(net127),
    .B1_N(net147),
    .X(net164));
 sky130_fd_sc_hd__a41o_1 c240 (.A1(net164),
    .A2(net151),
    .A3(net114),
    .A4(net882),
    .B1(net878),
    .X(net165));
 sky130_fd_sc_hd__a31o_1 c241 (.A1(net156),
    .A2(net882),
    .A3(net161),
    .B1(net676),
    .X(net166));
 sky130_fd_sc_hd__a21bo_1 c242 (.A1(net111),
    .A2(net32),
    .B1_N(net44),
    .X(net167));
 sky130_fd_sc_hd__a21bo_1 c243 (.A1(net159),
    .A2(net841),
    .B1_N(net896),
    .X(net168));
 sky130_fd_sc_hd__a41o_1 c244 (.A1(net148),
    .A2(net783),
    .A3(net882),
    .A4(net131),
    .B1(net32),
    .X(net169));
 sky130_fd_sc_hd__a21bo_2 c245 (.A1(net50),
    .A2(net779),
    .B1_N(net798),
    .X(net871));
 sky130_fd_sc_hd__a21bo_1 c246 (.A1(net42),
    .A2(net870),
    .B1_N(net32),
    .X(net170));
 sky130_fd_sc_hd__a41o_1 c247 (.A1(net818),
    .A2(net169),
    .A3(net135),
    .A4(net45),
    .B1(net871),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net32),
    .A1(net37),
    .A2(net126),
    .A3(net864),
    .S0(net863),
    .S1(net882),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net760),
    .X(net872));
 sky130_fd_sc_hd__a41o_1 c250 (.A1(net780),
    .A2(net811),
    .A3(net871),
    .A4(net872),
    .B1(net850),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 c251 (.A(net978),
    .X(net174));
 sky130_fd_sc_hd__sdfbbp_1 c252 (.CLK(clknet_4_5_0_clk),
    .D(net126),
    .RESET_B(net780),
    .SCD(net36),
    .SCE(net871),
    .SET_B(net163),
    .Q(net176),
    .Q_N(net175));
 sky130_fd_sc_hd__a41o_1 c253 (.A1(net168),
    .A2(net813),
    .A3(net866),
    .A4(net811),
    .B1(net830),
    .X(net177));
 sky130_fd_sc_hd__a21bo_1 c254 (.A1(net131),
    .A2(net50),
    .B1_N(net882),
    .X(net178));
 sky130_fd_sc_hd__a21bo_1 c255 (.A1(net791),
    .A2(net870),
    .B1_N(net148),
    .X(net179));
 sky130_fd_sc_hd__sdfbbn_1 c256 (.CLK_N(clknet_4_4_0_clk),
    .D(net179),
    .RESET_B(net171),
    .SCD(net45),
    .SCE(net783),
    .SET_B(net168),
    .Q(net848),
    .Q_N(net180));
 sky130_fd_sc_hd__a41o_1 c257 (.A1(net143),
    .A2(net848),
    .A3(net178),
    .A4(net163),
    .B1(net780),
    .X(net181));
 sky130_fd_sc_hd__a21bo_1 c258 (.A1(net176),
    .A2(net36),
    .B1_N(net37),
    .X(net844));
 sky130_fd_sc_hd__sdfbbn_1 c259 (.CLK_N(clknet_4_4_0_clk),
    .D(net174),
    .RESET_B(net173),
    .SCD(net871),
    .SCE(net844),
    .SET_B(net980),
    .Q(net868));
 sky130_fd_sc_hd__sdfbbp_1 c260 (.CLK(clknet_4_4_0_clk),
    .D(net44),
    .RESET_B(net122),
    .SCD(net178),
    .SCE(net635),
    .SET_B(net179),
    .Q(net842));
 sky130_fd_sc_hd__clkbuf_1 c261 (.A(net761),
    .X(net854));
 sky130_fd_sc_hd__a21bo_1 c262 (.A1(net871),
    .A2(net3),
    .B1_N(net658),
    .X(net182));
 sky130_fd_sc_hd__a41o_1 c263 (.A1(net122),
    .A2(net170),
    .A3(net866),
    .A4(net635),
    .B1(net175),
    .X(net183));
 sky130_fd_sc_hd__xnor2_2 c264 (.A(net777),
    .B(net915),
    .Y(net184));
 sky130_fd_sc_hd__xnor2_4 c265 (.A(net1000),
    .B(net832),
    .Y(net185));
 sky130_fd_sc_hd__a21bo_2 c266 (.A1(net769),
    .A2(net71),
    .B1_N(net185),
    .X(net186));
 sky130_fd_sc_hd__xnor2_4 c267 (.A(net63),
    .B(net902),
    .Y(net187));
 sky130_fd_sc_hd__xnor2_1 c268 (.A(net72),
    .B(net773),
    .Y(net857));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net187),
    .B(net73),
    .Y(net188));
 sky130_fd_sc_hd__xnor2_2 c270 (.A(net81),
    .B(net919),
    .Y(net189));
 sky130_fd_sc_hd__xnor2_4 c271 (.A(net913),
    .B(net906),
    .Y(net190));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net903),
    .B(net925),
    .Y(net191));
 sky130_fd_sc_hd__a41o_4 c273 (.A1(net190),
    .A2(net894),
    .A3(net78),
    .A4(net63),
    .B1(net902),
    .X(net192));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net895),
    .B(net906),
    .Y(net193));
 sky130_fd_sc_hd__xnor2_2 c275 (.A(net185),
    .B(net192),
    .Y(net194));
 sky130_fd_sc_hd__a21bo_4 c276 (.A1(net894),
    .A2(net194),
    .B1_N(net895),
    .X(net195));
 sky130_fd_sc_hd__a31o_4 c277 (.A1(net186),
    .A2(net1000),
    .A3(net190),
    .B1(net194),
    .X(net196));
 sky130_fd_sc_hd__xnor2_4 c278 (.A(net900),
    .B(net941),
    .Y(net837));
 sky130_fd_sc_hd__xnor2_4 c279 (.A(net195),
    .B(net193),
    .Y(net197));
 sky130_fd_sc_hd__a41o_4 c280 (.A1(net888),
    .A2(net837),
    .A3(net906),
    .A4(net196),
    .B1(net895),
    .X(net198));
 sky130_fd_sc_hd__xnor2_4 c281 (.A(net192),
    .B(net191),
    .Y(net199));
 sky130_fd_sc_hd__xnor2_2 c282 (.A(net900),
    .B(net888),
    .Y(net200));
 sky130_fd_sc_hd__xnor2_4 c283 (.A(net196),
    .B(net198),
    .Y(net201));
 sky130_fd_sc_hd__a41o_4 c284 (.A1(net201),
    .A2(net900),
    .A3(net772),
    .A4(net894),
    .B1(net915),
    .X(net853));
 sky130_fd_sc_hd__a31o_1 c285 (.A1(net73),
    .A2(net201),
    .A3(net907),
    .B1(net200),
    .X(net202));
 sky130_fd_sc_hd__xnor2_4 c286 (.A(net895),
    .B(net921),
    .Y(net203));
 sky130_fd_sc_hd__xnor2_4 c287 (.A(net960),
    .B(net796),
    .Y(net204));
 sky130_fd_sc_hd__a21bo_4 c288 (.A1(net203),
    .A2(net185),
    .B1_N(net921),
    .X(net205));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net202),
    .A2(net803),
    .B1_N(net906),
    .X(net860));
 sky130_fd_sc_hd__xnor2_4 c290 (.A(net780),
    .B(net203),
    .Y(net206));
 sky130_fd_sc_hd__xnor2_4 c291 (.A(net185),
    .B(net888),
    .Y(net207));
 sky130_fd_sc_hd__xnor2_1 c292 (.A(net206),
    .B(net97),
    .Y(net208));
 sky130_fd_sc_hd__xnor2_2 c293 (.A(net805),
    .B(net199),
    .Y(net209));
 sky130_fd_sc_hd__mux4_2 c294 (.A0(net775),
    .A1(net205),
    .A2(net93),
    .A3(net91),
    .S0(net207),
    .S1(net204),
    .X(net210));
 sky130_fd_sc_hd__xnor2_4 c295 (.A(net96),
    .B(net210),
    .Y(net211));
 sky130_fd_sc_hd__a41o_2 c296 (.A1(net80),
    .A2(net74),
    .A3(net204),
    .A4(net958),
    .B1(net921),
    .X(net212));
 sky130_fd_sc_hd__xnor2_4 c297 (.A(net942),
    .B(net205),
    .Y(net213));
 sky130_fd_sc_hd__xnor2_1 c298 (.A(net211),
    .B(net83),
    .Y(net214));
 sky130_fd_sc_hd__xnor2_4 c299 (.A(net213),
    .B(net211),
    .Y(net215));
 sky130_fd_sc_hd__a41o_2 c300 (.A1(net85),
    .A2(net215),
    .A3(net211),
    .A4(net209),
    .B1(net920),
    .X(net216));
 sky130_fd_sc_hd__a21bo_2 c301 (.A1(net215),
    .A2(net213),
    .B1_N(net205),
    .X(net217));
 sky130_fd_sc_hd__buf_2 c302 (.A(net763),
    .X(net218));
 sky130_fd_sc_hd__a31o_1 c303 (.A1(net209),
    .A2(net205),
    .A3(net860),
    .B1(net218),
    .X(net219));
 sky130_fd_sc_hd__a41o_1 c304 (.A1(net217),
    .A2(net204),
    .A3(net215),
    .A4(net198),
    .B1(net207),
    .X(net220));
 sky130_fd_sc_hd__a31o_1 c305 (.A1(net888),
    .A2(net208),
    .A3(net218),
    .B1(net895),
    .X(net221));
 sky130_fd_sc_hd__a21bo_1 c306 (.A1(net87),
    .A2(net221),
    .B1_N(net211),
    .X(net222));
 sky130_fd_sc_hd__a31o_1 c307 (.A1(net202),
    .A2(net860),
    .A3(net216),
    .B1(net219),
    .X(net223));
 sky130_fd_sc_hd__xnor2_1 c308 (.A(net821),
    .B(net652),
    .Y(net224));
 sky130_fd_sc_hd__a41o_2 c309 (.A1(net768),
    .A2(net219),
    .A3(net221),
    .A4(net779),
    .B1(net776),
    .X(net225));
 sky130_fd_sc_hd__a31o_1 c310 (.A1(net797),
    .A2(net204),
    .A3(net78),
    .B1(net207),
    .X(net226));
 sky130_fd_sc_hd__a21bo_4 c311 (.A1(net210),
    .A2(net1013),
    .B1_N(net997),
    .X(net227));
 sky130_fd_sc_hd__xnor2_2 c312 (.A(net998),
    .B(net799),
    .Y(net228));
 sky130_fd_sc_hd__xnor2_1 c313 (.A(net780),
    .B(net84),
    .Y(net229));
 sky130_fd_sc_hd__a21bo_1 c314 (.A1(net806),
    .A2(net91),
    .B1_N(net825),
    .X(net230));
 sky130_fd_sc_hd__xnor2_4 c315 (.A(net107),
    .B(net227),
    .Y(net231));
 sky130_fd_sc_hd__a21bo_2 c316 (.A1(net203),
    .A2(net228),
    .B1_N(net816),
    .X(net232));
 sky130_fd_sc_hd__a21bo_1 c317 (.A1(net84),
    .A2(net218),
    .B1_N(net224),
    .X(net233));
 sky130_fd_sc_hd__a21bo_4 c318 (.A1(net110),
    .A2(net958),
    .B1_N(net233),
    .X(net234));
 sky130_fd_sc_hd__a21bo_1 c319 (.A1(net219),
    .A2(net232),
    .B1_N(net652),
    .X(net235));
 sky130_fd_sc_hd__xnor2_1 c320 (.A(net209),
    .B(net772),
    .Y(net236));
 sky130_fd_sc_hd__xnor2_4 c321 (.A(net232),
    .B(net84),
    .Y(net237));
 sky130_fd_sc_hd__a21bo_1 c322 (.A1(net237),
    .A2(net203),
    .B1_N(net652),
    .X(net238));
 sky130_fd_sc_hd__buf_2 c323 (.A(net672),
    .X(net239));
 sky130_fd_sc_hd__xnor2_4 c324 (.A(net234),
    .B(net807),
    .Y(net852));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net238),
    .A1(net78),
    .A2(net226),
    .A3(net225),
    .S0(net915),
    .S1(net652),
    .X(net240));
 sky130_fd_sc_hd__a21bo_2 c326 (.A1(net226),
    .A2(net229),
    .B1_N(net677),
    .X(net241));
 sky130_fd_sc_hd__a41o_4 c327 (.A1(net109),
    .A2(net230),
    .A3(net238),
    .A4(net815),
    .B1(net228),
    .X(net855));
 sky130_fd_sc_hd__mux4_1 c328 (.A0(net236),
    .A1(net915),
    .A2(net241),
    .A3(net855),
    .S0(net234),
    .S1(net920),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net242),
    .A1(net1),
    .A2(net237),
    .A3(net234),
    .S0(net209),
    .S1(net225),
    .X(net243));
 sky130_fd_sc_hd__a31o_4 c330 (.A1(net184),
    .A2(net867),
    .A3(net104),
    .B1(net20),
    .X(net244));
 sky130_fd_sc_hd__a21bo_1 c331 (.A1(net959),
    .A2(net207),
    .B1_N(net19),
    .X(net245));
 sky130_fd_sc_hd__mux4_2 c332 (.A0(net120),
    .A1(net78),
    .A2(net234),
    .A3(net241),
    .S0(net900),
    .S1(net806),
    .X(net246));
 sky130_fd_sc_hd__sdfbbn_1 c333 (.CLK_N(clknet_4_0_0_clk),
    .D(net130),
    .RESET_B(net246),
    .SCD(net921),
    .SCE(net9),
    .SET_B(net883),
    .Q(net248),
    .Q_N(net247));
 sky130_fd_sc_hd__a31o_1 c334 (.A1(net244),
    .A2(net213),
    .A3(net864),
    .B1(net959),
    .X(net249));
 sky130_fd_sc_hd__sdfrbp_1 c335 (.CLK(clknet_4_0_0_clk),
    .D(net246),
    .RESET_B(net241),
    .SCD(net799),
    .SCE(net883),
    .Q(net251),
    .Q_N(net250));
 sky130_fd_sc_hd__sdfbbn_1 c336 (.CLK_N(clknet_4_0_0_clk),
    .D(net977),
    .RESET_B(net130),
    .SCD(net120),
    .SCE(net246),
    .SET_B(net816),
    .Q(net253),
    .Q_N(net252));
 sky130_fd_sc_hd__a41o_1 c337 (.A1(net241),
    .A2(net852),
    .A3(net82),
    .A4(net855),
    .B1(net247),
    .X(net254));
 sky130_fd_sc_hd__mux4_2 c338 (.A0(net249),
    .A1(net953),
    .A2(net137),
    .A3(net245),
    .S0(net892),
    .S1(net678),
    .X(net255));
 sky130_fd_sc_hd__a21bo_1 c339 (.A1(net224),
    .A2(net227),
    .B1_N(net252),
    .X(net256));
 sky130_fd_sc_hd__a21bo_1 c340 (.A1(net83),
    .A2(net860),
    .B1_N(net207),
    .X(net257));
 sky130_fd_sc_hd__a31o_1 c341 (.A1(net972),
    .A2(net257),
    .A3(net130),
    .B1(net988),
    .X(net258));
 sky130_fd_sc_hd__sdfbbp_1 c342 (.CLK(clknet_4_1_0_clk),
    .D(net256),
    .RESET_B(net972),
    .SCD(net118),
    .SCE(net883),
    .SET_B(net970),
    .Q(net260),
    .Q_N(net259));
 sky130_fd_sc_hd__sdfbbn_1 c343 (.CLK_N(clknet_4_1_0_clk),
    .D(net260),
    .RESET_B(net255),
    .SCD(net878),
    .SCE(net212),
    .SET_B(net1010),
    .Q(net875),
    .Q_N(net261));
 sky130_fd_sc_hd__a31o_1 c344 (.A1(net933),
    .A2(net249),
    .A3(net254),
    .B1(net678),
    .X(net262));
 sky130_fd_sc_hd__a31o_1 c345 (.A1(net253),
    .A2(net87),
    .A3(net135),
    .B1(net245),
    .X(net263));
 sky130_fd_sc_hd__a31o_1 c346 (.A1(net213),
    .A2(net248),
    .A3(net878),
    .B1(net234),
    .X(net264));
 sky130_fd_sc_hd__a31o_1 c347 (.A1(net78),
    .A2(net104),
    .A3(net135),
    .B1(net257),
    .X(net265));
 sky130_fd_sc_hd__a31o_1 c348 (.A1(net258),
    .A2(net782),
    .A3(net979),
    .B1(net265),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net254),
    .A1(net262),
    .A2(net922),
    .A3(net96),
    .S0(net258),
    .S1(net892),
    .X(net267));
 sky130_fd_sc_hd__sdfbbn_1 c350 (.CLK_N(clknet_4_1_0_clk),
    .D(net260),
    .RESET_B(net265),
    .SCD(net184),
    .SCE(net245),
    .SET_B(net973),
    .Q(net268));
 sky130_fd_sc_hd__sdfrbp_1 c351 (.CLK(clknet_4_0_0_clk),
    .D(net265),
    .RESET_B(net268),
    .SCD(net259),
    .SCE(net115),
    .Q(net270),
    .Q_N(net269));
 sky130_fd_sc_hd__mux4_2 c352 (.A0(net166),
    .A1(net768),
    .A2(net82),
    .A3(net821),
    .S0(net824),
    .S1(net922),
    .X(net271));
 sky130_fd_sc_hd__a41o_1 c353 (.A1(net114),
    .A2(net92),
    .A3(net31),
    .A4(net82),
    .B1(net136),
    .X(net272));
 sky130_fd_sc_hd__a21bo_1 c354 (.A1(net7),
    .A2(net38),
    .B1_N(net855),
    .X(net273));
 sky130_fd_sc_hd__a41o_1 c355 (.A1(net115),
    .A2(net930),
    .A3(net859),
    .A4(net954),
    .B1(net162),
    .X(net274));
 sky130_fd_sc_hd__a41o_1 c356 (.A1(net129),
    .A2(net922),
    .A3(net231),
    .A4(net273),
    .B1(net31),
    .X(net275));
 sky130_fd_sc_hd__buf_1 c357 (.A(net626),
    .X(net276));
 sky130_fd_sc_hd__a41o_1 c358 (.A1(net161),
    .A2(net244),
    .A3(net24),
    .A4(net125),
    .B1(net199),
    .X(net277));
 sky130_fd_sc_hd__sdfrtn_1 c359 (.CLK_N(clknet_4_1_0_clk),
    .D(net125),
    .RESET_B(net793),
    .SCD(net271),
    .SCE(net985),
    .Q(net278));
 sky130_fd_sc_hd__a31o_1 c360 (.A1(net272),
    .A2(net9),
    .A3(net798),
    .B1(net38),
    .X(net279));
 sky130_fd_sc_hd__sdfbbp_1 c361 (.CLK(clknet_4_5_0_clk),
    .D(net157),
    .RESET_B(net816),
    .SCD(net156),
    .SCE(net273),
    .SET_B(net891),
    .Q(net281),
    .Q_N(net280));
 sky130_fd_sc_hd__a31o_1 c362 (.A1(net137),
    .A2(net855),
    .A3(net852),
    .B1(net278),
    .X(net840));
 sky130_fd_sc_hd__a31o_1 c363 (.A1(net136),
    .A2(net7),
    .A3(net244),
    .B1(net80),
    .X(net282));
 sky130_fd_sc_hd__a41o_2 c364 (.A1(net92),
    .A2(net859),
    .A3(net75),
    .A4(net261),
    .B1(net840),
    .X(net283));
 sky130_fd_sc_hd__buf_1 c365 (.A(net625),
    .X(net846));
 sky130_fd_sc_hd__sdfbbn_1 c366 (.CLK_N(clknet_4_5_0_clk),
    .D(net113),
    .RESET_B(net23),
    .SCD(net7),
    .SCE(net891),
    .SET_B(net283),
    .Q(net285),
    .Q_N(net284));
 sky130_fd_sc_hd__sdfbbn_1 c367 (.CLK_N(clknet_4_5_0_clk),
    .D(net158),
    .RESET_B(net281),
    .SCD(net283),
    .SCE(net801),
    .SET_B(net166),
    .Q(net287),
    .Q_N(net286));
 sky130_fd_sc_hd__sdfbbp_1 c368 (.CLK(clknet_4_7_0_clk),
    .D(net801),
    .RESET_B(net113),
    .SCD(net191),
    .SCE(net283),
    .SET_B(net890),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__sdfbbn_1 c369 (.CLK_N(clknet_4_7_0_clk),
    .D(net82),
    .RESET_B(net262),
    .SCD(net859),
    .SCE(net784),
    .SET_B(net288),
    .Q(net291),
    .Q_N(net290));
 sky130_fd_sc_hd__a41o_1 c370 (.A1(net273),
    .A2(net824),
    .A3(net287),
    .A4(net290),
    .B1(net160),
    .X(net292));
 sky130_fd_sc_hd__sdfrtp_1 c371 (.CLK(clknet_4_5_0_clk),
    .D(net283),
    .RESET_B(net965),
    .SCD(net982),
    .SCE(net668),
    .Q(net293));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(net162),
    .A1(net291),
    .A2(net293),
    .A3(net840),
    .S0(net284),
    .S1(net288),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_1 c373 (.A(net761),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net819),
    .A1(net60),
    .A2(net178),
    .A3(net135),
    .S0(net896),
    .S1(net811),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net167),
    .A1(net49),
    .A2(net829),
    .A3(net289),
    .S0(net58),
    .S1(net663),
    .X(net861));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net56),
    .A1(net863),
    .A2(net58),
    .A3(net664),
    .S0(net674),
    .S1(net858),
    .X(net862));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net135),
    .A1(net182),
    .A2(net874),
    .A3(net819),
    .S0(net867),
    .S1(net658),
    .X(net869));
 sky130_fd_sc_hd__xnor2_2 c396 (.A(net190),
    .B(net81),
    .Y(net296));
 sky130_fd_sc_hd__a21bo_4 c397 (.A1(net827),
    .A2(net192),
    .B1_N(net187),
    .X(net297));
 sky130_fd_sc_hd__xnor2_2 c398 (.A(net790),
    .B(net894),
    .Y(net298));
 sky130_fd_sc_hd__a21bo_4 c399 (.A1(net66),
    .A2(net190),
    .B1_N(net297),
    .X(net299));
 sky130_fd_sc_hd__xnor2_4 c400 (.A(net936),
    .B(net80),
    .Y(net833));
 sky130_fd_sc_hd__xnor2_4 c401 (.A(net197),
    .B(net833),
    .Y(net300));
 sky130_fd_sc_hd__xnor2_2 c402 (.A(net297),
    .B(net298),
    .Y(net301));
 sky130_fd_sc_hd__xnor2_2 c403 (.A(net300),
    .B(net299),
    .Y(net302));
 sky130_fd_sc_hd__xnor2_4 c404 (.A(net828),
    .B(net913),
    .Y(net303));
 sky130_fd_sc_hd__a21bo_1 c405 (.A1(net303),
    .A2(net296),
    .B1_N(net884),
    .X(net304));
 sky130_fd_sc_hd__a21bo_4 c406 (.A1(net304),
    .A2(net71),
    .B1_N(net885),
    .X(net305));
 sky130_fd_sc_hd__a41o_1 c407 (.A1(net305),
    .A2(net297),
    .A3(net197),
    .A4(net195),
    .B1(net884),
    .X(net306));
 sky130_fd_sc_hd__a21bo_2 c408 (.A1(net776),
    .A2(net303),
    .B1_N(net884),
    .X(net307));
 sky130_fd_sc_hd__a21bo_2 c409 (.A1(net298),
    .A2(net307),
    .B1_N(net884),
    .X(net308));
 sky130_fd_sc_hd__xnor2_2 c410 (.A(net307),
    .B(net308),
    .Y(net309));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(net300),
    .A2(net308),
    .B1_N(net884),
    .X(net310));
 sky130_fd_sc_hd__a31o_1 c412 (.A1(net301),
    .A2(net310),
    .A3(net938),
    .B1(net884),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 c413 (.A(net647),
    .X(net312));
 sky130_fd_sc_hd__a21bo_1 c414 (.A1(net884),
    .A2(net306),
    .B1_N(net903),
    .X(net313));
 sky130_fd_sc_hd__sdfrtp_4 c415 (.CLK(clknet_4_8_0_clk),
    .D(net313),
    .RESET_B(net971),
    .SCD(net308),
    .SCE(net307),
    .Q(net314));
 sky130_fd_sc_hd__a41o_1 c416 (.A1(net309),
    .A2(net310),
    .A3(net967),
    .A4(net196),
    .B1(net313),
    .X(net315));
 sky130_fd_sc_hd__sdfbbn_2 c417 (.CLK_N(clknet_4_8_0_clk),
    .D(net314),
    .RESET_B(net313),
    .SCD(net312),
    .SCE(net884),
    .SET_B(net646),
    .Q(net317),
    .Q_N(net316));
 sky130_fd_sc_hd__xnor2_2 c418 (.A(net773),
    .B(net91),
    .Y(net318));
 sky130_fd_sc_hd__a21bo_4 c419 (.A1(net192),
    .A2(net989),
    .B1_N(net884),
    .X(net319));
 sky130_fd_sc_hd__a21bo_1 c420 (.A1(net309),
    .A2(net97),
    .B1_N(net88),
    .X(net320));
 sky130_fd_sc_hd__xnor2_4 c421 (.A(net853),
    .B(net319),
    .Y(net321));
 sky130_fd_sc_hd__a41o_1 c422 (.A1(net307),
    .A2(net316),
    .A3(net940),
    .A4(net303),
    .B1(net800),
    .X(net322));
 sky130_fd_sc_hd__buf_1 c423 (.A(net662),
    .X(net323));
 sky130_fd_sc_hd__xnor2_4 c424 (.A(net828),
    .B(net787),
    .Y(net324));
 sky130_fd_sc_hd__a31o_2 c425 (.A1(net800),
    .A2(net911),
    .A3(net768),
    .B1(net62),
    .X(net325));
 sky130_fd_sc_hd__a31o_2 c426 (.A1(net208),
    .A2(net222),
    .A3(net905),
    .B1(net911),
    .X(net326));
 sky130_fd_sc_hd__a21bo_2 c427 (.A1(net911),
    .A2(net794),
    .B1_N(net921),
    .X(net327));
 sky130_fd_sc_hd__a21bo_1 c428 (.A1(net905),
    .A2(net319),
    .B1_N(net221),
    .X(net328));
 sky130_fd_sc_hd__a41o_1 c429 (.A1(net214),
    .A2(net322),
    .A3(net62),
    .A4(net889),
    .B1(net69),
    .X(net329));
 sky130_fd_sc_hd__a31o_2 c430 (.A1(net64),
    .A2(net88),
    .A3(net796),
    .B1(net309),
    .X(net330));
 sky130_fd_sc_hd__a21bo_2 c431 (.A1(net327),
    .A2(net64),
    .B1_N(net911),
    .X(net331));
 sky130_fd_sc_hd__a41o_2 c432 (.A1(net331),
    .A2(net194),
    .A3(net80),
    .A4(net305),
    .B1(net323),
    .X(net332));
 sky130_fd_sc_hd__buf_6 c433 (.A(net661),
    .X(net333));
 sky130_fd_sc_hd__mux4_2 c434 (.A0(net187),
    .A1(net323),
    .A2(net796),
    .A3(net307),
    .S0(net905),
    .S1(net887),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(net329),
    .A1(net218),
    .A2(net332),
    .A3(net918),
    .S0(net787),
    .S1(net328),
    .X(net335));
 sky130_fd_sc_hd__a41o_1 c436 (.A1(net823),
    .A2(net328),
    .A3(net911),
    .A4(net334),
    .B1(net903),
    .X(net336));
 sky130_fd_sc_hd__mux4_2 c437 (.A0(net332),
    .A1(net904),
    .A2(net336),
    .A3(net952),
    .S0(net911),
    .S1(net680),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net330),
    .A1(net307),
    .A2(net905),
    .A3(net329),
    .S0(net90),
    .S1(net316),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net332),
    .A1(net328),
    .A2(net329),
    .A3(net337),
    .S0(net905),
    .S1(clknet_1_0__leaf_net681),
    .X(net339));
 sky130_fd_sc_hd__dlymetal6s2s_1 c440 (.A(net650),
    .X(net851));
 sky130_fd_sc_hd__a31o_1 c441 (.A1(net91),
    .A2(net241),
    .A3(net813),
    .B1(net770),
    .X(net340));
 sky130_fd_sc_hd__a21bo_1 c442 (.A1(net221),
    .A2(net961),
    .B1_N(net646),
    .X(net341));
 sky130_fd_sc_hd__a31o_1 c443 (.A1(net852),
    .A2(net233),
    .A3(net327),
    .B1(net673),
    .X(net342));
 sky130_fd_sc_hd__a41o_1 c444 (.A1(net323),
    .A2(net200),
    .A3(net317),
    .A4(net904),
    .B1(net222),
    .X(net343));
 sky130_fd_sc_hd__a21bo_1 c445 (.A1(net222),
    .A2(net961),
    .B1_N(net234),
    .X(net344));
 sky130_fd_sc_hd__a21bo_1 c446 (.A1(net233),
    .A2(net186),
    .B1_N(net940),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 c447 (.A(net650),
    .X(net346));
 sky130_fd_sc_hd__a21bo_4 c448 (.A1(net992),
    .A2(net908),
    .B1_N(net662),
    .X(net873));
 sky130_fd_sc_hd__a21bo_1 c449 (.A1(net342),
    .A2(net233),
    .B1_N(net795),
    .X(net347));
 sky130_fd_sc_hd__a21bo_1 c450 (.A1(net317),
    .A2(net212),
    .B1_N(net867),
    .X(net348));
 sky130_fd_sc_hd__a31o_1 c451 (.A1(net310),
    .A2(net314),
    .A3(net908),
    .B1(net652),
    .X(net349));
 sky130_fd_sc_hd__a31o_4 c452 (.A1(net229),
    .A2(net234),
    .A3(net873),
    .B1(net881),
    .X(net350));
 sky130_fd_sc_hd__sdfbbp_1 c453 (.CLK(clknet_4_9_0_clk),
    .D(net348),
    .RESET_B(net905),
    .SCD(net347),
    .SCE(net238),
    .SET_B(net855),
    .Q(net352),
    .Q_N(net351));
 sky130_fd_sc_hd__sdfbbn_1 c454 (.CLK_N(clknet_4_9_0_clk),
    .D(net349),
    .RESET_B(net887),
    .SCD(net196),
    .SCE(net881),
    .SET_B(net343),
    .Q(net354),
    .Q_N(net353));
 sky130_fd_sc_hd__a41o_1 c455 (.A1(net345),
    .A2(net809),
    .A3(net354),
    .A4(net350),
    .B1(net348),
    .X(net355));
 sky130_fd_sc_hd__a21bo_1 c456 (.A1(net200),
    .A2(net69),
    .B1_N(net241),
    .X(net356));
 sky130_fd_sc_hd__a31o_4 c457 (.A1(net346),
    .A2(net105),
    .A3(net887),
    .B1(net650),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net797),
    .A1(net343),
    .A2(net350),
    .A3(net357),
    .S0(net353),
    .S1(net650),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net343),
    .A1(net191),
    .A2(net357),
    .A3(net881),
    .S0(net921),
    .S1(clknet_1_0__leaf_net682),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net72),
    .A1(net350),
    .A2(net90),
    .A3(net239),
    .S0(net357),
    .S1(clknet_1_0__leaf_net682),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net347),
    .A1(net350),
    .A2(net306),
    .A3(net357),
    .S0(clknet_1_0__leaf_net682),
    .S1(net684),
    .X(net361));
 sky130_fd_sc_hd__a41o_1 c462 (.A1(net875),
    .A2(net883),
    .A3(net820),
    .A4(net635),
    .B1(net685),
    .X(net362));
 sky130_fd_sc_hd__a31o_1 c463 (.A1(net964),
    .A2(net350),
    .A3(net362),
    .B1(net881),
    .X(net363));
 sky130_fd_sc_hd__a41o_2 c464 (.A1(net322),
    .A2(net269),
    .A3(net112),
    .A4(net80),
    .B1(net921),
    .X(net364));
 sky130_fd_sc_hd__sdfbbn_1 c465 (.CLK_N(clknet_4_3_0_clk),
    .D(net344),
    .RESET_B(net96),
    .SCD(net20),
    .SCE(net261),
    .SET_B(net263),
    .Q(net366),
    .Q_N(net365));
 sky130_fd_sc_hd__sdfbbp_1 c466 (.CLK(clknet_4_3_0_clk),
    .D(net262),
    .RESET_B(net852),
    .SCD(net795),
    .SCE(net883),
    .SET_B(net687),
    .Q(net368),
    .Q_N(net367));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(net366),
    .A1(net948),
    .A2(net118),
    .A3(net943),
    .S0(net679),
    .S1(net685),
    .X(net369));
 sky130_fd_sc_hd__a41o_1 c468 (.A1(net72),
    .A2(net364),
    .A3(net88),
    .A4(net879),
    .B1(net649),
    .X(net370));
 sky130_fd_sc_hd__sdfbbn_1 c469 (.CLK_N(clknet_4_6_0_clk),
    .D(net370),
    .RESET_B(net6),
    .SCD(net891),
    .SCE(net357),
    .SET_B(net879),
    .Q(net372),
    .Q_N(net371));
 sky130_fd_sc_hd__a41o_1 c470 (.A1(net934),
    .A2(net367),
    .A3(net318),
    .A4(net199),
    .B1(net852),
    .X(net373));
 sky130_fd_sc_hd__a41o_1 c471 (.A1(net306),
    .A2(net781),
    .A3(net932),
    .A4(net879),
    .B1(net371),
    .X(net374));
 sky130_fd_sc_hd__a41o_1 c472 (.A1(net1012),
    .A2(net813),
    .A3(net883),
    .A4(net357),
    .B1(net879),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net19),
    .A1(net256),
    .A2(net364),
    .A3(net875),
    .S0(net356),
    .S1(net879),
    .X(net376));
 sky130_fd_sc_hd__a41o_1 c474 (.A1(net228),
    .A2(net368),
    .A3(net365),
    .A4(net16),
    .B1(net684),
    .X(net377));
 sky130_fd_sc_hd__sdfbbn_1 c475 (.CLK_N(clknet_4_3_0_clk),
    .D(net915),
    .RESET_B(net235),
    .SCD(net813),
    .SCE(net6),
    .SET_B(net879),
    .Q(net379),
    .Q_N(net378));
 sky130_fd_sc_hd__a41o_1 c476 (.A1(net375),
    .A2(net367),
    .A3(net879),
    .A4(net1),
    .B1(clknet_1_0__leaf_net682),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 c477 (.A0(net377),
    .A1(net379),
    .A2(net9),
    .A3(net799),
    .S0(net364),
    .S1(net879),
    .X(net381));
 sky130_fd_sc_hd__a41o_1 c478 (.A1(net20),
    .A2(net372),
    .A3(net199),
    .A4(net195),
    .B1(net908),
    .X(net382));
 sky130_fd_sc_hd__a41o_1 c479 (.A1(net96),
    .A2(net250),
    .A3(net1003),
    .A4(net378),
    .B1(net646),
    .X(net383));
 sky130_fd_sc_hd__mux4_2 c480 (.A0(net787),
    .A1(net356),
    .A2(net364),
    .A3(net881),
    .S0(net879),
    .S1(net648),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net368),
    .A1(net382),
    .A2(net326),
    .A3(net384),
    .S0(net381),
    .S1(net686),
    .X(net385));
 sky130_fd_sc_hd__sdfbbp_1 c482 (.CLK(clknet_4_6_0_clk),
    .D(net383),
    .RESET_B(net199),
    .SCD(net370),
    .SCE(net384),
    .SET_B(net690),
    .Q(net387),
    .Q_N(net386));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net245),
    .A1(net383),
    .A2(net375),
    .A3(net384),
    .S0(clknet_1_0__leaf_net681),
    .S1(net688),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net292),
    .A1(net72),
    .A2(net282),
    .A3(net271),
    .S0(net830),
    .S1(net769),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 c485 (.A0(net160),
    .A1(net232),
    .A2(net386),
    .A3(net827),
    .S0(net843),
    .S1(net72),
    .X(net390));
 sky130_fd_sc_hd__sdfbbn_1 c486 (.CLK_N(clknet_4_6_0_clk),
    .D(net156),
    .RESET_B(net856),
    .SCD(net80),
    .SCE(net289),
    .SET_B(net384),
    .Q(net392),
    .Q_N(net391));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net191),
    .A1(net317),
    .A2(net828),
    .A3(net276),
    .S0(net813),
    .S1(net292),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c488 (.A0(net283),
    .A1(net776),
    .A2(net274),
    .A3(net824),
    .S0(net88),
    .S1(clknet_1_1__leaf_net681),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net80),
    .A1(net987),
    .A2(net34),
    .A3(net393),
    .S0(net810),
    .S1(net680),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net821),
    .A1(net867),
    .A2(net882),
    .A3(net922),
    .S0(clknet_1_1__leaf_net681),
    .S1(net692),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net824),
    .A1(clknet_1_0__leaf_net396),
    .A2(net852),
    .A3(net922),
    .S0(net946),
    .S1(net834),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net354),
    .A1(net390),
    .A2(net846),
    .A3(net391),
    .S0(net150),
    .S1(net892),
    .X(net398));
 sky130_fd_sc_hd__a41o_1 c493 (.A1(net795),
    .A2(net830),
    .A3(net828),
    .A4(net945),
    .B1(net687),
    .X(net847));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net199),
    .A1(net392),
    .A2(net384),
    .A3(net833),
    .S0(net24),
    .S1(net881),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net397),
    .A1(net856),
    .A2(net867),
    .A3(net277),
    .S0(net890),
    .S1(net696),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net373),
    .A1(net207),
    .A2(net847),
    .A3(net294),
    .S0(net244),
    .S1(net691),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net134),
    .A1(net395),
    .A2(net232),
    .A3(net635),
    .S0(net288),
    .S1(net851),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net387),
    .A1(net271),
    .A2(net794),
    .A3(net160),
    .S0(net887),
    .S1(net847),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(net207),
    .A1(net294),
    .A2(net326),
    .A3(net289),
    .S0(net887),
    .S1(net882),
    .X(net403));
 sky130_fd_sc_hd__sdfbbn_1 c500 (.CLK_N(clknet_4_7_0_clk),
    .D(net326),
    .RESET_B(net784),
    .SCD(net783),
    .SCE(net384),
    .SET_B(net923),
    .Q(net404));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net31),
    .A1(net283),
    .A2(net947),
    .A3(net261),
    .S0(net691),
    .S1(net983),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c502 (.A0(net150),
    .A1(net373),
    .A2(net294),
    .A3(net911),
    .S0(net955),
    .S1(net674),
    .X(net406));
 sky130_fd_sc_hd__a41o_1 c503 (.A1(net833),
    .A2(net930),
    .A3(net288),
    .A4(net923),
    .B1(net657),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net384),
    .A1(net830),
    .A2(net271),
    .A3(net956),
    .S0(net647),
    .S1(net984),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(net407),
    .A1(net316),
    .A2(net836),
    .A3(net288),
    .S0(net697),
    .S1(net698),
    .X(net409));
 sky130_fd_sc_hd__xnor2_4 c528 (.A(net916),
    .B(net926),
    .Y(net410));
 sky130_fd_sc_hd__xnor2_4 c529 (.A(net312),
    .B(net299),
    .Y(net411));
 sky130_fd_sc_hd__xnor2_1 c530 (.A(net296),
    .B(net777),
    .Y(net412));
 sky130_fd_sc_hd__clkbuf_2 c531 (.X(net413));
 sky130_fd_sc_hd__clkbuf_2 c532 (.A(net636),
    .X(net414));
 sky130_fd_sc_hd__a21bo_1 c533 (.A1(net919),
    .A2(net1015),
    .B1_N(net777),
    .X(net415));
 sky130_fd_sc_hd__xnor2_4 c534 (.A(net635),
    .B(net910),
    .Y(net877));
 sky130_fd_sc_hd__a21bo_4 c535 (.A1(net298),
    .A2(net413),
    .B1_N(net894),
    .X(net831));
 sky130_fd_sc_hd__xnor2_4 c536 (.A(net877),
    .B(net410),
    .Y(net416));
 sky130_fd_sc_hd__xnor2_4 c537 (.A(net893),
    .B(net910),
    .Y(net417));
 sky130_fd_sc_hd__xnor2_4 c538 (.A(net823),
    .B(net776),
    .Y(net418));
 sky130_fd_sc_hd__xnor2_4 c539 (.A(net910),
    .B(net416),
    .Y(net419));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(net66),
    .A2(net303),
    .B1_N(net894),
    .X(net420));
 sky130_fd_sc_hd__xnor2_2 c541 (.A(net415),
    .B(net908),
    .Y(net421));
 sky130_fd_sc_hd__xnor2_4 c542 (.A(net299),
    .B(net297),
    .Y(net422));
 sky130_fd_sc_hd__a21bo_1 c543 (.A1(net301),
    .A2(net304),
    .B1_N(net416),
    .X(net423));
 sky130_fd_sc_hd__xnor2_4 c544 (.A(net770),
    .B(net831),
    .Y(net424));
 sky130_fd_sc_hd__a21bo_2 c545 (.A1(net420),
    .A2(net424),
    .B1_N(net416),
    .X(net425));
 sky130_fd_sc_hd__mux4_2 c546 (.A0(net424),
    .A1(net421),
    .A2(net423),
    .A3(net66),
    .S0(net416),
    .S1(net410),
    .X(net426));
 sky130_fd_sc_hd__mux4_2 c547 (.A0(net304),
    .A1(net296),
    .A2(net424),
    .A3(net423),
    .S0(net831),
    .S1(net417),
    .X(net427));
 sky130_fd_sc_hd__a21bo_1 c548 (.A1(net421),
    .A2(net832),
    .B1_N(net1016),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net427),
    .A1(net420),
    .A2(net424),
    .A3(net428),
    .S0(net418),
    .S1(net421),
    .X(net429));
 sky130_fd_sc_hd__dlymetal6s2s_1 c550 (.A(net759),
    .X(net430));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net430),
    .A2(net411),
    .B1_N(net918),
    .X(net431));
 sky130_fd_sc_hd__a21bo_1 c552 (.A1(net427),
    .A2(net910),
    .B1_N(net425),
    .X(net432));
 sky130_fd_sc_hd__xnor2_4 c553 (.A(net903),
    .B(net417),
    .Y(net433));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net794),
    .B(net950),
    .Y(net434));
 sky130_fd_sc_hd__a21bo_1 c555 (.A1(net336),
    .A2(net430),
    .B1_N(net416),
    .X(net435));
 sky130_fd_sc_hd__a21bo_1 c556 (.A1(net300),
    .A2(net308),
    .B1_N(net905),
    .X(net436));
 sky130_fd_sc_hd__a21bo_1 c557 (.A1(net416),
    .A2(net891),
    .B1_N(net436),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 c558 (.A(net759),
    .X(net438));
 sky130_fd_sc_hd__a41o_1 c559 (.A1(net438),
    .A2(net911),
    .A3(net430),
    .A4(net889),
    .B1(net1026),
    .X(net439));
 sky130_fd_sc_hd__buf_1 c560 (.A(net763),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 c561 (.A(net672),
    .X(net441));
 sky130_fd_sc_hd__a31o_1 c562 (.A1(net415),
    .A2(net205),
    .A3(net434),
    .B1(net905),
    .X(net442));
 sky130_fd_sc_hd__a41o_1 c563 (.A1(net431),
    .A2(net777),
    .A3(net986),
    .A4(net319),
    .B1(net418),
    .X(net443));
 sky130_fd_sc_hd__a21bo_1 c564 (.A1(net417),
    .A2(net430),
    .B1_N(net431),
    .X(net444));
 sky130_fd_sc_hd__buf_1 c565 (.A(net766),
    .X(net445));
 sky130_fd_sc_hd__a21bo_2 c566 (.A1(net440),
    .A2(net438),
    .B1_N(net445),
    .X(net446));
 sky130_fd_sc_hd__mux4_2 c567 (.A0(net439),
    .A1(net422),
    .A2(net899),
    .A3(net440),
    .S0(net212),
    .S1(net797),
    .X(net839));
 sky130_fd_sc_hd__sdfrtp_1 c568 (.CLK(clknet_4_8_0_clk),
    .D(net435),
    .RESET_B(net336),
    .SCD(net331),
    .SCE(net899),
    .Q(net447));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net441),
    .A1(net447),
    .A2(net437),
    .A3(net950),
    .S0(net779),
    .S1(net899),
    .X(net448));
 sky130_fd_sc_hd__a41o_1 c570 (.A1(net966),
    .A2(net303),
    .A3(net442),
    .A4(net433),
    .B1(net899),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net429),
    .A1(net337),
    .A2(net447),
    .A3(net336),
    .S0(net961),
    .S1(net899),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 c572 (.A(net669),
    .X(net451));
 sky130_fd_sc_hd__a21bo_2 c573 (.A1(net97),
    .A2(net412),
    .B1_N(net939),
    .X(net452));
 sky130_fd_sc_hd__a21bo_1 c574 (.A1(net318),
    .A2(net825),
    .B1_N(net651),
    .X(net453));
 sky130_fd_sc_hd__a21bo_1 c575 (.A1(net412),
    .A2(net797),
    .B1_N(net2),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 c576 (.A(net669),
    .X(net455));
 sky130_fd_sc_hd__a21bo_1 c577 (.A1(net352),
    .A2(net924),
    .B1_N(net912),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c578 (.A(net762),
    .X(net457));
 sky130_fd_sc_hd__a21bo_1 c579 (.A1(net410),
    .A2(net839),
    .B1_N(net773),
    .X(net458));
 sky130_fd_sc_hd__a41o_1 c580 (.A1(net809),
    .A2(net309),
    .A3(net451),
    .A4(net904),
    .B1(net425),
    .X(net459));
 sky130_fd_sc_hd__a21bo_1 c581 (.A1(net89),
    .A2(net196),
    .B1_N(net453),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 c582 (.A(net762),
    .X(net461));
 sky130_fd_sc_hd__a41o_1 c583 (.A1(net230),
    .A2(net195),
    .A3(net833),
    .A4(net805),
    .B1(clknet_1_0__leaf_net683),
    .X(net462));
 sky130_fd_sc_hd__a21bo_1 c584 (.A1(net196),
    .A2(net204),
    .B1_N(net899),
    .X(net463));
 sky130_fd_sc_hd__a31o_1 c585 (.A1(net116),
    .A2(net823),
    .A3(net452),
    .B1(net899),
    .X(net464));
 sky130_fd_sc_hd__a41o_1 c586 (.A1(net464),
    .A2(net424),
    .A3(net438),
    .A4(net461),
    .B1(net831),
    .X(net465));
 sky130_fd_sc_hd__a21bo_1 c587 (.A1(net460),
    .A2(net781),
    .B1_N(net204),
    .X(net466));
 sky130_fd_sc_hd__a41o_1 c588 (.A1(net436),
    .A2(net833),
    .A3(net205),
    .A4(net899),
    .B1(net700),
    .X(net467));
 sky130_fd_sc_hd__a21bo_1 c589 (.A1(net463),
    .A2(net2),
    .B1_N(net651),
    .X(net468));
 sky130_fd_sc_hd__a41o_1 c590 (.A1(net899),
    .A2(net460),
    .A3(net904),
    .A4(net352),
    .B1(clknet_1_0__leaf_net462),
    .X(net469));
 sky130_fd_sc_hd__a21bo_1 c591 (.A1(net319),
    .A2(net799),
    .B1_N(net881),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net453),
    .A1(net990),
    .A2(net452),
    .A3(clknet_1_0__leaf_net469),
    .S0(net351),
    .S1(net470),
    .X(net471));
 sky130_fd_sc_hd__a41o_1 c593 (.A1(net461),
    .A2(net465),
    .A3(net468),
    .A4(net776),
    .B1(net899),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net467),
    .A1(clknet_1_0__leaf_net462),
    .A2(net422),
    .A3(net112),
    .S0(net364),
    .S1(net836),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net443),
    .A1(net991),
    .A2(net949),
    .A3(net1002),
    .S0(net892),
    .S1(net880),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net16),
    .A1(net816),
    .A2(net467),
    .A3(net1005),
    .S0(net939),
    .S1(net690),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net205),
    .A1(net374),
    .A2(net816),
    .A3(net112),
    .S0(net924),
    .S1(clknet_1_0__leaf_net701),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net827),
    .A1(net474),
    .A2(net426),
    .A3(net963),
    .S0(clknet_1_0__leaf_net683),
    .S1(clknet_1_1__leaf_net701),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net948),
    .A1(net889),
    .A2(net318),
    .A3(net16),
    .S0(net689),
    .S1(clknet_1_0__leaf_net702),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net458),
    .A1(net112),
    .A2(net893),
    .A3(net451),
    .S0(net820),
    .S1(clknet_1_1__leaf_net702),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net212),
    .A1(net244),
    .A2(net324),
    .A3(net234),
    .S0(net1001),
    .S1(clknet_1_0__leaf_net702),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net356),
    .A1(net479),
    .A2(net452),
    .A3(clknet_1_0__leaf_net480),
    .S0(net470),
    .S1(clknet_1_0__leaf_net702),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net270),
    .A1(net374),
    .A2(clknet_1_0__leaf_net478),
    .A3(net878),
    .S0(net770),
    .S1(net775),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net297),
    .A1(net1),
    .A2(net206),
    .A3(net878),
    .S0(net883),
    .S1(clknet_1_0__leaf_net478),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net112),
    .A1(net362),
    .A2(net794),
    .A3(net364),
    .S0(net18),
    .S1(clknet_1_0__leaf_net702),
    .X(net484));
 sky130_fd_sc_hd__mux4_2 c606 (.A0(net815),
    .A1(net836),
    .A2(net775),
    .A3(net880),
    .S0(net919),
    .S1(clknet_1_0__leaf_net682),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net71),
    .A1(clknet_1_1__leaf_net462),
    .A2(net795),
    .A3(net827),
    .S0(net667),
    .S1(clknet_1_0__leaf_net702),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net426),
    .A1(clknet_1_1__leaf_net480),
    .A2(clknet_1_0__leaf_net485),
    .A3(net889),
    .S0(net873),
    .S1(clknet_1_1__leaf_net702),
    .X(net487));
 sky130_fd_sc_hd__mux4_2 c609 (.A0(net321),
    .A1(clknet_1_1__leaf_net478),
    .A2(net795),
    .A3(net451),
    .S0(net893),
    .S1(clknet_1_1__leaf_net702),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net924),
    .A1(net486),
    .A2(net16),
    .A3(net422),
    .S0(net944),
    .S1(net635),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net364),
    .A1(clknet_1_1__leaf_net485),
    .A2(net451),
    .A3(net883),
    .S0(clknet_1_1__leaf_net702),
    .S1(net706),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net318),
    .A1(net470),
    .A2(net426),
    .A3(net350),
    .S0(net422),
    .S1(net364),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net910),
    .A1(net769),
    .A2(net883),
    .A3(clknet_1_0__leaf_net485),
    .S0(net667),
    .S1(clknet_1_1__leaf_net702),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net775),
    .A1(net484),
    .A2(net910),
    .A3(net792),
    .S0(net790),
    .S1(clknet_1_0__leaf_net702),
    .X(net492));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(net488),
    .A1(net771),
    .A2(net16),
    .A3(net990),
    .S0(clknet_1_1__leaf_net702),
    .S1(net710),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net24),
    .A1(net770),
    .A2(net400),
    .A3(net908),
    .S0(net779),
    .S1(net878),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(net350),
    .A1(net407),
    .A2(net945),
    .A3(net263),
    .S0(net919),
    .S1(net911),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net293),
    .A1(net18),
    .A2(net779),
    .A3(net879),
    .S0(net881),
    .S1(net669),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net423),
    .A1(net466),
    .A2(net404),
    .A3(net231),
    .S0(net890),
    .S1(net969),
    .X(net497));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net808),
    .A1(net786),
    .A2(net810),
    .A3(net824),
    .S0(net2),
    .S1(net818),
    .X(net0));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net425),
    .A1(net75),
    .A2(net793),
    .A3(net289),
    .S0(net768),
    .S1(net830),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net393),
    .A1(net9),
    .A2(clknet_1_1__leaf_net396),
    .A3(net892),
    .S0(net890),
    .S1(net878),
    .X(net499));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(net419),
    .A1(net11),
    .A2(net498),
    .A3(net88),
    .S0(net18),
    .S1(net873),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net878),
    .A1(net195),
    .A2(net880),
    .A3(net419),
    .S0(net11),
    .S1(net656),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net102),
    .A1(net468),
    .A2(net882),
    .A3(net836),
    .S0(net444),
    .S1(net711),
    .X(net502));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(net149),
    .A1(net263),
    .A2(net195),
    .A3(net793),
    .S0(net206),
    .S1(net838),
    .X(net503));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(net289),
    .A1(net794),
    .A2(net500),
    .A3(net836),
    .S0(net878),
    .S1(net882),
    .X(net504));
 sky130_fd_sc_hd__mux4_2 c627 (.A0(net218),
    .A1(net155),
    .A2(net890),
    .A3(net88),
    .S0(net878),
    .S1(net9),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net496),
    .A1(net880),
    .A2(net918),
    .A3(net770),
    .S0(net890),
    .S1(net357),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net276),
    .A1(net769),
    .A2(net890),
    .A3(net71),
    .S0(net798),
    .S1(net882),
    .X(net507));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net817),
    .A1(net821),
    .A2(net806),
    .A3(net816),
    .S0(net824),
    .S1(net818),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net444),
    .A1(net451),
    .A2(net195),
    .A3(net144),
    .S0(net75),
    .S1(net24),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net277),
    .A1(net1005),
    .A2(net24),
    .A3(net880),
    .S0(net770),
    .S1(net707),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net88),
    .A1(net771),
    .A2(net144),
    .A3(net880),
    .S0(net11),
    .S1(net703),
    .X(net510));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net425),
    .A1(net244),
    .A2(net880),
    .A3(net693),
    .S0(net714),
    .S1(net718),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net502),
    .A1(net472),
    .A2(net635),
    .A3(net289),
    .S0(net799),
    .S1(net700),
    .X(net512));
 sky130_fd_sc_hd__mux4_2 c635 (.A0(net507),
    .A1(net106),
    .A2(net498),
    .A3(net2),
    .S0(net793),
    .S1(net714),
    .X(net513));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net509),
    .A1(net324),
    .A2(net106),
    .A3(net350),
    .S0(net679),
    .S1(net711),
    .X(net514));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net278),
    .A1(net409),
    .A2(net830),
    .A3(net834),
    .S0(net716),
    .S1(net720),
    .X(net515));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net803),
    .A1(net819),
    .A2(net800),
    .A3(net815),
    .S0(net816),
    .S1(net820),
    .X(net1));
 sky130_fd_sc_hd__a41o_4 c65 (.A1(net785),
    .A2(net789),
    .A3(net774),
    .A4(net782),
    .B1(net798),
    .X(net2));
 sky130_fd_sc_hd__xnor2_2 c66 (.A(net787),
    .B(net810),
    .Y(net3));
 sky130_fd_sc_hd__a21bo_1 c660 (.A1(net777),
    .A2(net305),
    .B1_N(net411),
    .X(net516));
 sky130_fd_sc_hd__xnor2_4 c661 (.A(net812),
    .B(net305),
    .Y(net517));
 sky130_fd_sc_hd__xnor2_1 c662 (.A(net1018),
    .B(net908),
    .Y(net518));
 sky130_fd_sc_hd__a21bo_1 c663 (.A1(net790),
    .A2(net1017),
    .B1_N(net428),
    .X(net519));
 sky130_fd_sc_hd__xnor2_4 c664 (.A(net1024),
    .B(net81),
    .Y(net520));
 sky130_fd_sc_hd__a21bo_1 c665 (.A1(net516),
    .A2(net422),
    .B1_N(net424),
    .X(net521));
 sky130_fd_sc_hd__xnor2_1 c666 (.A(net428),
    .B(net771),
    .Y(net522));
 sky130_fd_sc_hd__buf_1 c667 (.A(net633),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_2 c668 (.A(net633),
    .X(net524));
 sky130_fd_sc_hd__a31o_1 c669 (.A1(net516),
    .A2(net907),
    .A3(net73),
    .B1(net1027),
    .X(net525));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net807),
    .B(net2),
    .Y(net4));
 sky130_fd_sc_hd__buf_1 c670 (.A(net665),
    .X(net526));
 sky130_fd_sc_hd__a21bo_1 c671 (.A1(net520),
    .A2(net517),
    .B1_N(net301),
    .X(net527));
 sky130_fd_sc_hd__xnor2_4 c672 (.A(net524),
    .B(net520),
    .Y(net528));
 sky130_fd_sc_hd__xnor2_2 c673 (.A(net414),
    .B(net528),
    .Y(net529));
 sky130_fd_sc_hd__clkbuf_1 c674 (.A(net665),
    .X(net530));
 sky130_fd_sc_hd__buf_2 c675 (.A(net647),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 c676 (.A(net765),
    .X(net532));
 sky130_fd_sc_hd__a21bo_1 c677 (.A1(net532),
    .A2(net427),
    .B1_N(net529),
    .X(net533));
 sky130_fd_sc_hd__a21bo_1 c678 (.A1(net529),
    .A2(net532),
    .B1_N(net530),
    .X(net534));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net528),
    .A1(net419),
    .A2(net532),
    .A3(net534),
    .S0(net912),
    .S1(net519),
    .X(net535));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net919),
    .B(net801),
    .Y(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 c680 (.A(net764),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(net534),
    .A1(net414),
    .A2(net533),
    .A3(net531),
    .S0(net532),
    .S1(net666),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 c682 (.A(net628),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net538),
    .A1(net189),
    .A2(net788),
    .A3(net217),
    .S0(net411),
    .S1(net680),
    .X(net539));
 sky130_fd_sc_hd__a21bo_1 c684 (.A1(net434),
    .A2(net1025),
    .B1_N(net834),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_1 c685 (.A(net627),
    .X(net541));
 sky130_fd_sc_hd__a21bo_1 c686 (.A1(net445),
    .A2(net517),
    .B1_N(net800),
    .X(net542));
 sky130_fd_sc_hd__a21bo_1 c687 (.A1(net526),
    .A2(net777),
    .B1_N(net433),
    .X(net543));
 sky130_fd_sc_hd__a21bo_1 c688 (.A1(net543),
    .A2(net186),
    .B1_N(net433),
    .X(net544));
 sky130_fd_sc_hd__sdfbbp_1 c689 (.CLK(clknet_4_8_0_clk),
    .D(net523),
    .RESET_B(net540),
    .SCD(net919),
    .SCE(net889),
    .SET_B(net898),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__xnor2_4 c69 (.A(net775),
    .B(net811),
    .Y(net864));
 sky130_fd_sc_hd__a31o_1 c690 (.A1(net518),
    .A2(net907),
    .A3(net898),
    .B1(net544),
    .X(net547));
 sky130_fd_sc_hd__sdfsbp_1 c691 (.CLK(clknet_4_10_0_clk),
    .D(net216),
    .SCD(net768),
    .SCE(net1027),
    .SET_B(net898),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__mux4_2 c692 (.A0(net902),
    .A1(net887),
    .A2(net518),
    .A3(net305),
    .S0(net308),
    .S1(net446),
    .X(net550));
 sky130_fd_sc_hd__a21bo_1 c693 (.A1(net541),
    .A2(net447),
    .B1_N(net331),
    .X(net551));
 sky130_fd_sc_hd__a41o_1 c694 (.A1(net951),
    .A2(net540),
    .A3(net420),
    .A4(net898),
    .B1(net542),
    .X(net552));
 sky130_fd_sc_hd__a21bo_1 c695 (.A1(net898),
    .A2(net531),
    .B1_N(net655),
    .X(net553));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net420),
    .A1(net331),
    .A2(net536),
    .A3(net433),
    .S0(net526),
    .S1(net332),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(net781),
    .A1(net216),
    .A2(net521),
    .A3(net189),
    .S0(net540),
    .S1(net553),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net554),
    .A1(net422),
    .A2(net327),
    .A3(net905),
    .S0(net721),
    .S1(net723),
    .X(net556));
 sky130_fd_sc_hd__mux4_2 c699 (.A0(net418),
    .A1(net427),
    .A2(net905),
    .A3(net327),
    .S0(net723),
    .S1(net725),
    .X(net557));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net5),
    .B(net787),
    .Y(net6));
 sky130_fd_sc_hd__a41o_2 c700 (.A1(net553),
    .A2(net548),
    .A3(net543),
    .A4(net898),
    .B1(net544),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net542),
    .A1(net414),
    .A2(net557),
    .A3(net543),
    .S0(net433),
    .S1(net554),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(net525),
    .A1(net434),
    .A2(net523),
    .A3(net558),
    .S0(net834),
    .S1(net726),
    .X(net560));
 sky130_fd_sc_hd__sdfbbn_1 c703 (.CLK_N(clknet_4_10_0_clk),
    .D(net549),
    .RESET_B(net445),
    .SCD(net558),
    .SCE(net557),
    .SET_B(net974),
    .Q(net562),
    .Q_N(net561));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net308),
    .A1(net330),
    .A2(net927),
    .A3(net204),
    .S0(net528),
    .S1(net887),
    .X(net563));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net800),
    .A1(net822),
    .A2(net898),
    .A3(net916),
    .S0(net1027),
    .S1(net330),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net557),
    .A1(net325),
    .A2(net771),
    .A3(net531),
    .S0(net545),
    .S1(net974),
    .X(net565));
 sky130_fd_sc_hd__mux4_2 c707 (.A0(net105),
    .A1(net516),
    .A2(net186),
    .A3(net418),
    .S0(net790),
    .S1(net550),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net531),
    .A1(net332),
    .A2(net820),
    .A3(net231),
    .S0(net889),
    .S1(net544),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net528),
    .A1(net546),
    .A2(net566),
    .A3(net898),
    .S0(clknet_1_1__leaf_net682),
    .S1(net727),
    .X(net568));
 sky130_fd_sc_hd__a21bo_1 c71 (.A1(net5),
    .A2(net768),
    .B1_N(net816),
    .X(net7));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net238),
    .A1(net424),
    .A2(net186),
    .A3(net517),
    .S0(net781),
    .S1(clknet_1_1__leaf_net683),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net411),
    .A1(net327),
    .A2(net557),
    .A3(net531),
    .S0(net536),
    .S1(net1028),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net465),
    .A1(net204),
    .A2(net822),
    .A3(net771),
    .S0(net652),
    .S1(net722),
    .X(net571));
 sky130_fd_sc_hd__mux4_2 c713 (.A0(net796),
    .A1(net215),
    .A2(net314),
    .A3(net544),
    .S0(net962),
    .S1(net728),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net805),
    .A1(net898),
    .A2(net419),
    .A3(net433),
    .S0(net561),
    .S1(net459),
    .X(net573));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net303),
    .A1(net798),
    .A2(net770),
    .A3(clknet_1_0__leaf_net469),
    .S0(net891),
    .S1(net186),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net433),
    .A1(net73),
    .A2(net572),
    .A3(net798),
    .S0(net545),
    .S1(net733),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net571),
    .A1(net797),
    .A2(net239),
    .A3(net452),
    .S0(net547),
    .S1(net446),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net777),
    .A1(net891),
    .A2(net807),
    .A3(net516),
    .S0(net727),
    .S1(net733),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net807),
    .A1(net419),
    .A2(net551),
    .A3(net733),
    .S0(net734),
    .S1(net735),
    .X(net578));
 sky130_fd_sc_hd__xnor2_1 c72 (.A(net806),
    .B(net6),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(net217),
    .A1(net825),
    .A2(net330),
    .A3(net898),
    .S0(net732),
    .S1(net734),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(net305),
    .A1(net577),
    .A2(net533),
    .A3(net908),
    .S0(net733),
    .S1(clknet_1_0__leaf_net736),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net237),
    .A1(net571),
    .A2(net889),
    .A3(net670),
    .S0(net733),
    .S1(clknet_1_1__leaf_net737),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net822),
    .A1(net578),
    .A2(net566),
    .A3(net531),
    .S0(net325),
    .S1(net733),
    .X(net582));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net544),
    .A1(clknet_1_0__leaf_net574),
    .A2(net61),
    .A3(net558),
    .S0(net724),
    .S1(net738),
    .X(net583));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net825),
    .A1(net583),
    .A2(net547),
    .A3(net225),
    .S0(clknet_1_0__leaf_net736),
    .S1(clknet_1_0__leaf_net737),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net540),
    .A1(net381),
    .A2(net790),
    .A3(net255),
    .S0(net546),
    .S1(net517),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net517),
    .A1(net769),
    .A2(net891),
    .A3(net709),
    .S0(net724),
    .S1(net742),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net533),
    .A1(net784),
    .A2(net776),
    .A3(net799),
    .S0(net708),
    .S1(net741),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net912),
    .A1(net255),
    .A2(net418),
    .A3(net438),
    .S0(net781),
    .S1(net700),
    .X(net588));
 sky130_fd_sc_hd__a21bo_4 c73 (.A1(net789),
    .A2(net864),
    .B1_N(net818),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net919),
    .A1(net381),
    .A2(net961),
    .A3(net891),
    .S0(net781),
    .S1(net722),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net820),
    .A1(net456),
    .A2(net929),
    .A3(net381),
    .S0(net919),
    .S1(net968),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net418),
    .A1(net186),
    .A2(net234),
    .A3(net781),
    .S0(clknet_1_1__leaf_net682),
    .S1(net729),
    .X(net591));
 sky130_fd_sc_hd__mux4_2 c733 (.A0(net904),
    .A1(net887),
    .A2(net808),
    .A3(clknet_1_1__leaf_net682),
    .S0(clknet_1_0__leaf_net737),
    .S1(net744),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net452),
    .A1(net784),
    .A2(net807),
    .A3(net680),
    .S0(clknet_1_1__leaf_net682),
    .S1(net733),
    .X(net593));
 sky130_fd_sc_hd__mux4_2 c735 (.A0(net883),
    .A1(net781),
    .A2(clknet_1_0__leaf_net592),
    .A3(net768),
    .S0(net653),
    .S1(net680),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net422),
    .A1(net536),
    .A2(clknet_1_1__leaf_net592),
    .A3(net558),
    .S0(net908),
    .S1(net788),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net551),
    .A1(net572),
    .A2(clknet_1_1__leaf_net469),
    .A3(net889),
    .S0(net690),
    .S1(net728),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net204),
    .A1(clknet_1_0__leaf_net592),
    .A2(clknet_1_0__leaf_net594),
    .A3(net572),
    .S0(net456),
    .S1(net726),
    .X(net597));
 sky130_fd_sc_hd__mux4_2 c739 (.A0(net547),
    .A1(net100),
    .A2(net773),
    .A3(clknet_1_1__leaf_net594),
    .S0(net781),
    .S1(clknet_1_1__leaf_net682),
    .X(net598));
 sky130_fd_sc_hd__a21bo_2 c74 (.A1(net864),
    .A2(net820),
    .B1_N(net6),
    .X(net10));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net455),
    .A1(net562),
    .A2(net142),
    .A3(net962),
    .S0(net726),
    .S1(net743),
    .X(net599));
 sky130_fd_sc_hd__mux4_2 c741 (.A0(net598),
    .A1(net928),
    .A2(net790),
    .A3(clknet_1_1__leaf_net469),
    .S0(net881),
    .S1(net743),
    .X(net600));
 sky130_fd_sc_hd__mux4_2 c742 (.A0(net225),
    .A1(net569),
    .A2(net314),
    .A3(clknet_1_0__leaf_net493),
    .S0(net419),
    .S1(net239),
    .X(net601));
 sky130_fd_sc_hd__mux4_2 c743 (.A0(net591),
    .A1(clknet_1_0__leaf_net600),
    .A2(net961),
    .A3(net517),
    .S0(net381),
    .S1(net690),
    .X(net602));
 sky130_fd_sc_hd__mux4_2 c744 (.A0(net550),
    .A1(net881),
    .A2(clknet_1_1__leaf_net600),
    .A3(net239),
    .S0(net654),
    .S1(net748),
    .X(net603));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net459),
    .A1(net808),
    .A2(clknet_1_0__leaf_net574),
    .A3(net768),
    .S0(net769),
    .S1(net741),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net227),
    .A1(net239),
    .A2(net79),
    .A3(net558),
    .S0(net709),
    .S1(net730),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net916),
    .A1(net225),
    .A2(net18),
    .A3(net726),
    .S0(net742),
    .S1(net976),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net457),
    .A1(net438),
    .A2(net795),
    .A3(net769),
    .S0(clknet_1_1__leaf_net683),
    .S1(clknet_1_1__leaf_net702),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(net595),
    .A1(net285),
    .A2(net103),
    .A3(net357),
    .S0(net694),
    .S1(net745),
    .X(net608));
 sky130_fd_sc_hd__xnor2_4 c75 (.A(net815),
    .B(net923),
    .Y(net11));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net558),
    .A1(net768),
    .A2(net902),
    .A3(net656),
    .S0(net692),
    .S1(net750),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net887),
    .A1(net593),
    .A2(net776),
    .A3(net607),
    .S0(net653),
    .S1(net705),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net788),
    .A1(net566),
    .A2(net799),
    .A3(net699),
    .S0(clknet_1_1__leaf_net719),
    .S1(net728),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net282),
    .A1(net918),
    .A2(net2),
    .A3(net896),
    .S0(net712),
    .S1(clknet_1_1__leaf_net736),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net546),
    .A1(net771),
    .A2(net788),
    .A3(net500),
    .S0(net752),
    .S1(net753),
    .X(net613));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net892),
    .A1(net274),
    .A2(clknet_1_1__leaf_net493),
    .A3(net771),
    .S0(net902),
    .S1(net739),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net340),
    .A1(net908),
    .A2(net206),
    .A3(net511),
    .S0(net613),
    .S1(net717),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net771),
    .A1(net911),
    .A2(net503),
    .A3(net744),
    .S0(net746),
    .S1(net755),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(net609),
    .A1(net34),
    .A2(net605),
    .A3(net599),
    .S0(net704),
    .S1(net731),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(net784),
    .A1(net810),
    .A2(clknet_1_1__leaf_net574),
    .A3(net608),
    .S0(net616),
    .S1(net700),
    .X(net618));
 sky130_fd_sc_hd__xnor2_2 c76 (.A(net6),
    .B(net776),
    .Y(net12));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net513),
    .A1(net239),
    .A2(clknet_1_1__leaf_net469),
    .A3(net610),
    .S0(clknet_1_0__leaf_net719),
    .S1(net749),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net357),
    .A1(net231),
    .A2(net896),
    .A3(net513),
    .S0(net715),
    .S1(net740),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net586),
    .A1(net79),
    .A2(net944),
    .A3(net515),
    .S0(net734),
    .S1(net757),
    .X(net621));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net799),
    .A1(net618),
    .A2(net680),
    .A3(net751),
    .S0(net756),
    .S1(net758),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net1005),
    .A1(net234),
    .A2(net619),
    .A3(net670),
    .S0(net713),
    .S1(net754),
    .X(net623));
 sky130_fd_sc_hd__a31o_2 c77 (.A1(net801),
    .A2(net0),
    .A3(net922),
    .B1(net10),
    .X(net13));
 sky130_fd_sc_hd__xnor2_4 c78 (.A(net804),
    .B(net897),
    .Y(net14));
 sky130_fd_sc_hd__a31o_4 c79 (.A1(net13),
    .A2(net6),
    .A3(net897),
    .B1(net922),
    .X(net15));
 sky130_fd_sc_hd__xnor2_2 c80 (.A(net1),
    .B(net4),
    .Y(net16));
 sky130_fd_sc_hd__xnor2_4 c81 (.A(net11),
    .B(net13),
    .Y(net17));
 sky130_fd_sc_hd__a41o_4 c82 (.A1(net897),
    .A2(net924),
    .A3(net836),
    .A4(net810),
    .B1(net804),
    .X(net843));
 sky130_fd_sc_hd__xnor2_4 c83 (.A(net17),
    .B(net14),
    .Y(net18));
 sky130_fd_sc_hd__a41o_2 c84 (.A1(net843),
    .A2(net1),
    .A3(net13),
    .A4(net0),
    .B1(net806),
    .X(net19));
 sky130_fd_sc_hd__a31o_2 c85 (.A1(net15),
    .A2(net785),
    .A3(net17),
    .B1(net922),
    .X(net856));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net6),
    .A1(net897),
    .A2(net15),
    .A3(net815),
    .S0(net19),
    .S1(net828),
    .X(net866));
 sky130_fd_sc_hd__a41o_2 c87 (.A1(net4),
    .A2(net11),
    .A3(net856),
    .A4(net866),
    .B1(net15),
    .X(net20));
 sky130_fd_sc_hd__xnor2_1 c88 (.A(net778),
    .B(net892),
    .Y(net21));
 sky130_fd_sc_hd__xnor2_4 c89 (.A(net772),
    .B(net9),
    .Y(net22));
 sky130_fd_sc_hd__a21bo_2 c90 (.A1(net4),
    .A2(net897),
    .B1_N(net21),
    .X(net23));
 sky130_fd_sc_hd__xnor2_4 c91 (.A(net798),
    .B(net772),
    .Y(net24));
 sky130_fd_sc_hd__a21bo_4 c92 (.A1(net21),
    .A2(net817),
    .B1_N(net816),
    .X(net830));
 sky130_fd_sc_hd__xnor2_4 c93 (.A(net23),
    .B(net15),
    .Y(net829));
 sky130_fd_sc_hd__a21bo_1 c94 (.A1(net22),
    .A2(net801),
    .B1_N(net830),
    .X(net25));
 sky130_fd_sc_hd__xnor2_4 c95 (.A(net15),
    .B(net4),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_1 c96 (.A(net779),
    .B(net26),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_4 c97 (.A(net26),
    .B(net782),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_4 c98 (.A(net829),
    .B(net28),
    .Y(net29));
 sky130_fd_sc_hd__xnor2_1 c99 (.A(net635),
    .B(net897),
    .Y(net30));
 sky130_fd_sc_hd__mux4_1 merge765 (.A0(net986),
    .A1(net429),
    .A2(net300),
    .A3(net437),
    .S0(net805),
    .S1(net1004),
    .X(net624));
 sky130_fd_sc_hd__sdfbbn_1 merge766 (.CLK_N(clknet_4_1_0_clk),
    .D(net257),
    .RESET_B(net246),
    .SCD(net772),
    .SCE(net773),
    .SET_B(net975),
    .Q(net626),
    .Q_N(net625));
 sky130_fd_sc_hd__sdfbbp_1 merge767 (.CLK(clknet_4_10_0_clk),
    .D(net521),
    .RESET_B(net517),
    .SCD(net419),
    .SCE(net894),
    .SET_B(net777),
    .Q(net628),
    .Q_N(net627));
 sky130_fd_sc_hd__mux4_1 merge768 (.A0(net320),
    .A1(net204),
    .A2(net235),
    .A3(net823),
    .S0(net652),
    .S1(net673),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 merge769 (.A0(net442),
    .A1(net112),
    .A2(net341),
    .A3(net89),
    .S0(net330),
    .S1(net652),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 merge770 (.A0(net146),
    .A1(net40),
    .A2(net147),
    .A3(net782),
    .S0(net122),
    .S1(net32),
    .X(net631));
 sky130_fd_sc_hd__a41o_1 merge771 (.A1(net795),
    .A2(net320),
    .A3(net322),
    .A4(net194),
    .B1(net912),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_1 merge772 (.A(net767),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 merge773 (.A0(net45),
    .A1(net172),
    .A2(net811),
    .A3(net57),
    .S0(net826),
    .S1(net49),
    .X(net634));
 sky130_fd_sc_hd__sdfbbn_2 merge774 (.CLK_N(clknet_4_8_0_clk),
    .D(net313),
    .SCD(net779),
    .SCE(net311),
    .SET_B(net1015),
    .Q(net636),
    .Q_N(net413));
 sky130_fd_sc_hd__a41o_1 merge775 (.A1(net525),
    .A2(net524),
    .A3(net528),
    .A4(net527),
    .B1(net523),
    .X(net637));
 sky130_fd_sc_hd__a41o_1 merge776 (.A1(net46),
    .A2(net53),
    .A3(net139),
    .A4(net113),
    .B1(net143),
    .X(net638));
 sky130_fd_sc_hd__mux4_1 merge777 (.A0(net311),
    .A1(net828),
    .A2(net884),
    .A3(net527),
    .S0(net529),
    .S1(net520),
    .X(net639));
 sky130_fd_sc_hd__mux4_1 merge778 (.A0(net280),
    .A1(net286),
    .A2(net865),
    .A3(net163),
    .S0(net37),
    .S1(net844),
    .X(net640));
 sky130_fd_sc_hd__mux4_1 merge779 (.A0(net90),
    .A1(net411),
    .A2(net442),
    .A3(net454),
    .S0(net350),
    .S1(net651),
    .X(net641));
 sky130_fd_sc_hd__mux4_1 merge780 (.A0(net331),
    .A1(net337),
    .A2(net334),
    .A3(net214),
    .S0(net216),
    .S1(net217),
    .X(net642));
 sky130_fd_sc_hd__mux4_1 merge781 (.A0(net121),
    .A1(net236),
    .A2(net902),
    .A3(net328),
    .S0(net435),
    .S1(net823),
    .X(net643));
 sky130_fd_sc_hd__mux4_1 merge782 (.A0(net530),
    .A1(net528),
    .A2(net525),
    .A3(net311),
    .S0(net532),
    .S1(net981),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 merge783 (.A0(net519),
    .A1(net522),
    .A2(net770),
    .A3(net432),
    .S0(net332),
    .S1(net438),
    .X(net645));
 sky130_fd_sc_hd__dfrbp_2 merge784 (.CLK(clknet_4_8_0_clk),
    .D(net639),
    .RESET_B(net315),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__dfrbp_1 merge785 (.CLK(clknet_4_3_0_clk),
    .D(net363),
    .RESET_B(net380),
    .Q(net649),
    .Q_N(net648));
 sky130_fd_sc_hd__dfrtn_1 merge786 (.CLK_N(clknet_4_2_0_clk),
    .D(net355),
    .RESET_B(net629),
    .Q(net650));
 sky130_fd_sc_hd__dfrtp_1 merge787 (.CLK(clknet_4_8_0_clk),
    .D(net448),
    .RESET_B(net449),
    .Q(net651));
 sky130_fd_sc_hd__dfrtp_1 merge788 (.CLK(clknet_4_0_0_clk),
    .RESET_B(net123),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 merge789 (.CLK(clknet_4_11_0_clk),
    .D(net589),
    .RESET_B(net590),
    .Q(net653));
 sky130_fd_sc_hd__dfsbp_1 merge790 (.CLK(clknet_4_14_0_clk),
    .D(net622),
    .SET_B(net623));
 sky130_fd_sc_hd__dfsbp_1 merge791 (.CLK(clknet_4_10_0_clk),
    .D(net539),
    .SET_B(net552),
    .Q(net655),
    .Q_N(net654));
 sky130_fd_sc_hd__dfstp_1 merge792 (.CLK(clknet_4_12_0_clk),
    .D(net494),
    .SET_B(net497),
    .Q(net656));
 sky130_fd_sc_hd__dfstp_1 merge793 (.CLK(clknet_4_7_0_clk),
    .D(net401),
    .SET_B(net402),
    .Q(net657));
 sky130_fd_sc_hd__dfstp_1 merge794 (.CLK(clknet_4_4_0_clk),
    .D(net177),
    .SET_B(net181),
    .Q(net658));
 sky130_fd_sc_hd__dlrbn_1 merge795 (.D(net165),
    .GATE_N(clknet_4_4_0_clk),
    .RESET_B(net631),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__dlrbn_1 merge796 (.D(net339),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net632),
    .Q(net662),
    .Q_N(net661));
 sky130_fd_sc_hd__dlrbp_1 merge797 (.D(net279),
    .GATE(clknet_4_5_0_clk),
    .RESET_B(net275),
    .Q(net664),
    .Q_N(net663));
 sky130_fd_sc_hd__dlrbp_1 merge798 (.D(net535),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net637),
    .Q(net666),
    .Q_N(net665));
 sky130_fd_sc_hd__dlrtn_1 merge799 (.D(net475),
    .GATE_N(clknet_4_12_0_clk),
    .RESET_B(net476),
    .Q(net667));
 sky130_fd_sc_hd__dlrtn_1 merge800 (.D(net264),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net266),
    .Q(net668));
 sky130_fd_sc_hd__dlrtn_1 merge801 (.D(net471),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net630),
    .Q(net669));
 sky130_fd_sc_hd__dlrtp_1 merge802 (.D(net563),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net564),
    .Q(net670));
 sky130_fd_sc_hd__dlrtp_1 merge803 (.D(net55),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net638),
    .Q(net671));
 sky130_fd_sc_hd__dlrtp_4 merge804 (.D(net223),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net220),
    .Q(net834));
 sky130_fd_sc_hd__edfxbp_1 merge805 (.CLK(clknet_4_2_0_clk),
    .D(net243),
    .DE(net643),
    .Q(net673),
    .Q_N(net672));
 sky130_fd_sc_hd__edfxtp_1 merge806 (.CLK(clknet_4_7_0_clk),
    .D(net403),
    .DE(net183),
    .Q(net674));
 sky130_fd_sc_hd__dfxbp_1 s807 (.CLK(clknet_4_4_0_clk),
    .D(net145),
    .Q(net676),
    .Q_N(net675));
 sky130_fd_sc_hd__dfxbp_1 s808 (.CLK(clknet_4_3_0_clk),
    .D(net240),
    .Q(net678),
    .Q_N(net677));
 sky130_fd_sc_hd__dfxtp_1 s809 (.CLK(clknet_4_1_0_clk),
    .D(net267),
    .Q(net679));
 sky130_fd_sc_hd__dfxtp_1 s810 (.CLK(clknet_4_5_0_clk),
    .D(net295),
    .Q(net858));
 sky130_fd_sc_hd__dfxtp_4 s811 (.CLK(clknet_4_2_0_clk),
    .D(net335),
    .Q(net680));
 sky130_fd_sc_hd__dlclkp_1 s812 (.CLK(clknet_4_2_0_clk),
    .GATE(net338),
    .GCLK(net681));
 sky130_fd_sc_hd__dlclkp_2 s813 (.CLK(clknet_4_9_0_clk),
    .GATE(net358),
    .GCLK(net682));
 sky130_fd_sc_hd__dlclkp_4 s814 (.CLK(clknet_4_9_0_clk),
    .GATE(net359),
    .GCLK(net683));
 sky130_fd_sc_hd__dlxbn_1 s815 (.D(net360),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__dlxbn_1 s816 (.D(net361),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__dlxbp_1 s817 (.D(net376),
    .GATE(clknet_4_3_0_clk),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dlxtn_2 s818 (.D(net385),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net690));
 sky130_fd_sc_hd__dlxtn_1 s819 (.D(net388),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net691));
 sky130_fd_sc_hd__dlxtn_1 s820 (.D(net389),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net692));
 sky130_fd_sc_hd__dlxtp_1 s821 (.D(net394),
    .GATE(clknet_4_7_0_clk),
    .Q(net693));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s822 (.D(net398),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net694));
 sky130_fd_sc_hd__dfxbp_1 s823 (.CLK(clknet_4_6_0_clk),
    .D(net399),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__dfxbp_1 s824 (.CLK(clknet_4_7_0_clk),
    .D(net405),
    .Q(net697));
 sky130_fd_sc_hd__dfxtp_1 s825 (.CLK(clknet_4_7_0_clk),
    .D(net406),
    .Q(net698));
 sky130_fd_sc_hd__dfxtp_1 s826 (.CLK(clknet_4_15_0_clk),
    .D(net408),
    .Q(net699));
 sky130_fd_sc_hd__dfxtp_2 s827 (.CLK(clknet_4_8_0_clk),
    .D(net450),
    .Q(net700));
 sky130_fd_sc_hd__dlclkp_1 s828 (.CLK(clknet_4_12_0_clk),
    .GATE(net473),
    .GCLK(net701));
 sky130_fd_sc_hd__dlclkp_2 s829 (.CLK(clknet_4_12_0_clk),
    .GATE(net477),
    .GCLK(net702));
 sky130_fd_sc_hd__dlclkp_4 s830 (.CLK(clknet_4_13_0_clk),
    .GATE(net481),
    .GCLK(net703));
 sky130_fd_sc_hd__dlxbn_1 s831 (.D(net482),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net876));
 sky130_fd_sc_hd__dlxbn_1 s832 (.D(net483),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net705),
    .Q_N(net704));
 sky130_fd_sc_hd__dlxbp_1 s833 (.D(net487),
    .GATE(clknet_4_12_0_clk),
    .Q(net707),
    .Q_N(net706));
 sky130_fd_sc_hd__dlxtn_1 s834 (.D(net489),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net708));
 sky130_fd_sc_hd__dlxtn_1 s835 (.D(net490),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net709));
 sky130_fd_sc_hd__dlxtn_1 s836 (.D(net491),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net710));
 sky130_fd_sc_hd__dlxtp_1 s837 (.D(net492),
    .GATE(clknet_4_6_0_clk),
    .Q(net838));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s838 (.D(net495),
    .SLEEP_B(clknet_4_13_0_clk),
    .Q(net711));
 sky130_fd_sc_hd__dfxbp_1 s839 (.CLK(clknet_4_13_0_clk),
    .D(net499),
    .Q(net712));
 sky130_fd_sc_hd__dfxbp_1 s840 (.CLK(clknet_4_15_0_clk),
    .D(net501),
    .Q(net713));
 sky130_fd_sc_hd__dfxtp_1 s841 (.CLK(clknet_4_13_0_clk),
    .D(net504),
    .Q(net714));
 sky130_fd_sc_hd__dfxtp_1 s842 (.CLK(clknet_4_15_0_clk),
    .D(net505),
    .Q(net715));
 sky130_fd_sc_hd__dfxtp_1 s843 (.CLK(clknet_4_13_0_clk),
    .D(net506),
    .Q(net716));
 sky130_fd_sc_hd__dlclkp_1 s844 (.CLK(clknet_4_13_0_clk),
    .GATE(net508),
    .GCLK(net717));
 sky130_fd_sc_hd__dlclkp_2 s845 (.CLK(clknet_4_13_0_clk),
    .GATE(net510),
    .GCLK(net718));
 sky130_fd_sc_hd__dlclkp_4 s846 (.CLK(clknet_4_15_0_clk),
    .GATE(net512),
    .GCLK(net719));
 sky130_fd_sc_hd__dlxbn_1 s847 (.D(net514),
    .GATE_N(clknet_4_13_0_clk),
    .Q(net720));
 sky130_fd_sc_hd__dlxbn_1 s848 (.D(net537),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net722),
    .Q_N(net721));
 sky130_fd_sc_hd__dlxbp_1 s849 (.D(net555),
    .GATE(clknet_4_10_0_clk),
    .Q(net724),
    .Q_N(net723));
 sky130_fd_sc_hd__dlxtn_1 s850 (.D(net556),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net725));
 sky130_fd_sc_hd__dlxtn_2 s851 (.D(net559),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net726));
 sky130_fd_sc_hd__dlxtn_1 s852 (.D(net560),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net727));
 sky130_fd_sc_hd__dlxtp_1 s853 (.D(net565),
    .GATE(clknet_4_10_0_clk),
    .Q(net728));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s854 (.D(net567),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net729));
 sky130_fd_sc_hd__dfxbp_1 s855 (.CLK(clknet_4_14_0_clk),
    .D(net568),
    .Q(net731),
    .Q_N(net730));
 sky130_fd_sc_hd__dfxbp_1 s856 (.CLK(clknet_4_10_0_clk),
    .D(net570),
    .Q(net732));
 sky130_fd_sc_hd__dfxtp_2 s857 (.CLK(clknet_4_10_0_clk),
    .D(net573),
    .Q(net733));
 sky130_fd_sc_hd__dfxtp_1 s858 (.CLK(clknet_4_11_0_clk),
    .D(net575),
    .Q(net734));
 sky130_fd_sc_hd__dfxtp_1 s859 (.CLK(clknet_4_11_0_clk),
    .D(net576),
    .Q(net735));
 sky130_fd_sc_hd__dlclkp_1 s860 (.CLK(clknet_4_11_0_clk),
    .GATE(net579),
    .GCLK(net736));
 sky130_fd_sc_hd__dlclkp_2 s861 (.CLK(clknet_4_11_0_clk),
    .GATE(net580),
    .GCLK(net737));
 sky130_fd_sc_hd__dlclkp_4 s862 (.CLK(clknet_4_11_0_clk),
    .GATE(net581),
    .GCLK(net738));
 sky130_fd_sc_hd__dlxbn_1 s863 (.D(net582),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net739));
 sky130_fd_sc_hd__dlxbn_1 s864 (.D(net584),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net740));
 sky130_fd_sc_hd__dlxbp_1 s865 (.D(net585),
    .GATE(clknet_4_14_0_clk),
    .Q(net742),
    .Q_N(net741));
 sky130_fd_sc_hd__dlxtn_1 s866 (.D(net587),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxtn_1 s867 (.D(net588),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net744));
 sky130_fd_sc_hd__dlxtn_1 s868 (.D(net596),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net745));
 sky130_fd_sc_hd__dlxtp_1 s869 (.D(net597),
    .GATE(clknet_4_15_0_clk),
    .Q(net746));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s870 (.D(net601),
    .SLEEP_B(clknet_4_14_0_clk),
    .Q(net747));
 sky130_fd_sc_hd__dfxbp_1 s871 (.CLK(clknet_4_11_0_clk),
    .D(net602),
    .Q(net748));
 sky130_fd_sc_hd__dfxbp_1 s872 (.CLK(clknet_4_14_0_clk),
    .D(net603),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_1 s873 (.CLK(clknet_4_12_0_clk),
    .D(net604),
    .Q(net750));
 sky130_fd_sc_hd__dfxtp_1 s874 (.CLK(clknet_4_14_0_clk),
    .D(net606),
    .Q(net751));
 sky130_fd_sc_hd__dfxtp_1 s875 (.CLK(clknet_4_15_0_clk),
    .D(net611),
    .Q(net752));
 sky130_fd_sc_hd__dlclkp_1 s876 (.CLK(clknet_4_13_0_clk),
    .GATE(net612),
    .GCLK(net753));
 sky130_fd_sc_hd__dlclkp_2 s877 (.CLK(clknet_4_14_0_clk),
    .GATE(net614),
    .GCLK(net754));
 sky130_fd_sc_hd__dlclkp_4 s878 (.CLK(clknet_4_13_0_clk),
    .GATE(net615),
    .GCLK(net755));
 sky130_fd_sc_hd__dlxbn_1 s879 (.D(net617),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net756));
 sky130_fd_sc_hd__dlxbn_1 s880 (.D(net620),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net757));
 sky130_fd_sc_hd__dlxbp_1 s881 (.D(net621),
    .GATE(clknet_4_15_0_clk),
    .Q(net758));
 sky130_fd_sc_hd__dlxtn_1 s882 (.D(net624),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net759));
 sky130_fd_sc_hd__dlxtn_1 s883 (.D(net634),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net760));
 sky130_fd_sc_hd__dlxtn_1 s884 (.D(net640),
    .GATE_N(clknet_4_7_0_clk),
    .Q(net761));
 sky130_fd_sc_hd__dlxtp_1 s885 (.D(net641),
    .GATE(clknet_4_9_0_clk),
    .Q(net762));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s886 (.D(net642),
    .SLEEP_B(clknet_4_8_0_clk),
    .Q(net763));
 sky130_fd_sc_hd__dfxbp_1 s887 (.CLK(clknet_4_10_0_clk),
    .D(net644),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dfxbp_1 s888 (.CLK(clknet_4_8_0_clk),
    .D(net645),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(in0),
    .X(net635));
 sky130_fd_sc_hd__buf_6 input2 (.A(in1),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(in10),
    .X(net769));
 sky130_fd_sc_hd__buf_12 input4 (.A(in11),
    .X(net770));
 sky130_fd_sc_hd__buf_4 input5 (.A(in12),
    .X(net771));
 sky130_fd_sc_hd__buf_8 input6 (.A(in13),
    .X(net772));
 sky130_fd_sc_hd__buf_12 input7 (.A(in14),
    .X(net773));
 sky130_fd_sc_hd__buf_6 input8 (.A(in15),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(in16),
    .X(net775));
 sky130_fd_sc_hd__buf_6 input10 (.A(in17),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(in18),
    .X(net777));
 sky130_fd_sc_hd__buf_8 input12 (.A(in19),
    .X(net778));
 sky130_fd_sc_hd__buf_4 input13 (.A(in2),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(in20),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(in21),
    .X(net781));
 sky130_fd_sc_hd__buf_4 input16 (.A(in22),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(in23),
    .X(net783));
 sky130_fd_sc_hd__buf_2 input18 (.A(in24),
    .X(net784));
 sky130_fd_sc_hd__buf_2 input19 (.A(in25),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_8 input21 (.A(in27),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(in28),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in29),
    .X(net789));
 sky130_fd_sc_hd__buf_12 input24 (.A(in3),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in30),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net793));
 sky130_fd_sc_hd__buf_2 input28 (.A(in33),
    .X(net794));
 sky130_fd_sc_hd__buf_4 input29 (.A(in34),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in35),
    .X(net796));
 sky130_fd_sc_hd__buf_2 input31 (.A(in36),
    .X(net797));
 sky130_fd_sc_hd__buf_6 input32 (.A(in37),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_8 input33 (.A(in38),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(in39),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(in4),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in40),
    .X(net802));
 sky130_fd_sc_hd__buf_2 input37 (.A(in41),
    .X(net803));
 sky130_fd_sc_hd__buf_4 input38 (.A(in42),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(in43),
    .X(net805));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net806));
 sky130_fd_sc_hd__buf_4 input41 (.A(in45),
    .X(net807));
 sky130_fd_sc_hd__buf_2 input42 (.A(in46),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in47),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(in48),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(in49),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_16 input46 (.A(in5),
    .X(net812));
 sky130_fd_sc_hd__buf_2 input47 (.A(in50),
    .X(net813));
 sky130_fd_sc_hd__buf_1 input48 (.A(in51),
    .X(net814));
 sky130_fd_sc_hd__buf_4 input49 (.A(in52),
    .X(net815));
 sky130_fd_sc_hd__buf_4 input50 (.A(in53),
    .X(net816));
 sky130_fd_sc_hd__buf_2 input51 (.A(in54),
    .X(net817));
 sky130_fd_sc_hd__buf_2 input52 (.A(in55),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in56),
    .X(net819));
 sky130_fd_sc_hd__buf_4 input54 (.A(in57),
    .X(net820));
 sky130_fd_sc_hd__buf_2 input55 (.A(in58),
    .X(net821));
 sky130_fd_sc_hd__buf_2 input56 (.A(in59),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(in6),
    .X(net823));
 sky130_fd_sc_hd__buf_2 input58 (.A(in60),
    .X(net824));
 sky130_fd_sc_hd__buf_2 input59 (.A(in61),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in7),
    .X(net826));
 sky130_fd_sc_hd__buf_6 input61 (.A(in8),
    .X(net827));
 sky130_fd_sc_hd__buf_6 input62 (.A(in9),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net829),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net830),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output65 (.A(net831),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output66 (.A(net896),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net833),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output68 (.A(net834),
    .X(out17));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net835),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net836),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output71 (.A(net993),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net838),
    .X(out20));
 sky130_fd_sc_hd__buf_2 output73 (.A(net839),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net840),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output75 (.A(net841),
    .X(out25));
 sky130_fd_sc_hd__buf_2 output76 (.A(net842),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output77 (.A(net843),
    .X(out28));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net844),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net845),
    .X(out3));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net846),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net847),
    .X(out31));
 sky130_fd_sc_hd__buf_2 output82 (.A(net848),
    .X(out32));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net849),
    .X(out33));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net850),
    .X(out35));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net851),
    .X(out36));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net852),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net955),
    .X(out38));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net854),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net855),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net856),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output91 (.A(net857),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net858),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net859),
    .X(out46));
 sky130_fd_sc_hd__buf_2 output94 (.A(net860),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net861),
    .X(out48));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net862),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output97 (.A(net863),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output98 (.A(net864),
    .X(out50));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net865),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net866),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output101 (.A(net867),
    .X(out53));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net868),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output103 (.A(net869),
    .X(out55));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net870),
    .X(out56));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net871),
    .X(out57));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net872),
    .X(out59));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net873),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output108 (.A(net874),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net875),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output110 (.A(net876),
    .X(out7));
 sky130_fd_sc_hd__buf_2 output111 (.A(net877),
    .X(out9));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(net144),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net369),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net369),
    .X(net880));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net340),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net835),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net142),
    .X(net883));
 sky130_fd_sc_hd__buf_12 fanout118 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__buf_12 fanout119 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(net302),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(net103),
    .X(net887));
 sky130_fd_sc_hd__buf_6 max_cap122 (.A(net197),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net100),
    .X(net889));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net106),
    .X(net890));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net102),
    .X(net891));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net18),
    .X(net892));
 sky130_fd_sc_hd__buf_4 max_cap127 (.A(net191),
    .X(net893));
 sky130_fd_sc_hd__buf_6 max_cap128 (.A(net189),
    .X(net894));
 sky130_fd_sc_hd__buf_12 fanout129 (.A(net188),
    .X(net895));
 sky130_fd_sc_hd__buf_4 wire130 (.A(net832),
    .X(net896));
 sky130_fd_sc_hd__buf_4 max_cap131 (.A(net12),
    .X(net897));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net446),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net446),
    .X(net899));
 sky130_fd_sc_hd__buf_4 max_cap134 (.A(net857),
    .X(net900));
 sky130_fd_sc_hd__buf_4 max_cap135 (.A(net82),
    .X(net901));
 sky130_fd_sc_hd__buf_12 max_cap136 (.A(net76),
    .X(net902));
 sky130_fd_sc_hd__buf_4 wire137 (.A(net74),
    .X(net903));
 sky130_fd_sc_hd__buf_8 fanout138 (.A(net333),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net325),
    .X(net905));
 sky130_fd_sc_hd__buf_4 max_cap140 (.A(net184),
    .X(net906));
 sky130_fd_sc_hd__buf_4 wire141 (.A(net79),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net68),
    .X(net908));
 sky130_fd_sc_hd__buf_6 max_cap143 (.A(net65),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_8 max_cap144 (.A(net413),
    .X(net910));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net324),
    .X(net911));
 sky130_fd_sc_hd__buf_6 max_cap146 (.A(net70),
    .X(net912));
 sky130_fd_sc_hd__buf_4 max_cap147 (.A(net936),
    .X(net913));
 sky130_fd_sc_hd__buf_6 max_cap148 (.A(net64),
    .X(net914));
 sky130_fd_sc_hd__buf_12 max_cap149 (.A(net63),
    .X(net915));
 sky130_fd_sc_hd__buf_6 max_cap150 (.A(net62),
    .X(net916));
 sky130_fd_sc_hd__buf_6 max_cap151 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_12 wire152 (.A(net61),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout153 (.A(net826),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net923),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net802),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net792),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net737 (.A(net737),
    .X(clknet_0_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_0__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net737 (.A(clknet_0_net737),
    .X(clknet_1_1__leaf_net737));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net592 (.A(net592),
    .X(clknet_0_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_0__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net592 (.A(clknet_0_net592),
    .X(clknet_1_1__leaf_net592));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net594 (.A(net594),
    .X(clknet_0_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_0__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net594 (.A(clknet_0_net594),
    .X(clknet_1_1__leaf_net594));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net736 (.A(net736),
    .X(clknet_0_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_0__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net736 (.A(clknet_0_net736),
    .X(clknet_1_1__leaf_net736));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net719 (.A(net719),
    .X(clknet_0_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_0__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net719 (.A(clknet_0_net719),
    .X(clknet_1_1__leaf_net719));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net480 (.A(net480),
    .X(clknet_0_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net480 (.A(clknet_0_net480),
    .X(clknet_1_0__leaf_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net480 (.A(clknet_0_net480),
    .X(clknet_1_1__leaf_net480));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net478 (.A(net478),
    .X(clknet_0_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_0__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net478 (.A(clknet_0_net478),
    .X(clknet_1_1__leaf_net478));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net701 (.A(net701),
    .X(clknet_0_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_0__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net701 (.A(clknet_0_net701),
    .X(clknet_1_1__leaf_net701));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net683 (.A(net683),
    .X(clknet_0_net683));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net683 (.A(clknet_0_net683),
    .X(clknet_1_0__leaf_net683));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net683 (.A(clknet_0_net683),
    .X(clknet_1_1__leaf_net683));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net462 (.A(net462),
    .X(clknet_0_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_0__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net462 (.A(clknet_0_net462),
    .X(clknet_1_1__leaf_net462));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net682 (.A(net682),
    .X(clknet_0_net682));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net682 (.A(clknet_0_net682),
    .X(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net682 (.A(clknet_0_net682),
    .X(clknet_1_1__leaf_net682));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net485 (.A(net485),
    .X(clknet_0_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_0__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net485 (.A(clknet_0_net485),
    .X(clknet_1_1__leaf_net485));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net681 (.A(net681),
    .X(clknet_0_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net681 (.A(clknet_0_net681),
    .X(clknet_1_1__leaf_net681));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net187),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net81),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net926),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net927),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net928),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net76),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net930),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer8 (.A(net935),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer9 (.A(net69),
    .X(net933));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer10 (.A(net933),
    .X(net934));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer11 (.A(net933),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net67),
    .X(net936));
 sky130_fd_sc_hd__buf_2 rebuffer13 (.A(net936),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net940),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer15 (.A(net940),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(net188),
    .X(net940));
 sky130_fd_sc_hd__buf_2 rebuffer17 (.A(net193),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net941),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net886),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net943),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net943),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net945),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net946),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(net188),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net948),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net334),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net950),
    .X(net951));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer28 (.A(net334),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net853),
    .X(net953));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer30 (.A(net953),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(net954),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(net955),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net70),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net198),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net958),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net198),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net962),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net333),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net337),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net963),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net288),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net447),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net314),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net733),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net694),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net834),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net312),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net251),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net668),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net726),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net660),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net747),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net248),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net760),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net259),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net180),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net666),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net664),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net695),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net693),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net660),
    .X(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A4 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_Y (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B1_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_Y (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_S0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_B1_N (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A4 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_A4 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_D (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_Y (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_SCE (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SET_B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCD (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_B1_N (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SCD (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_RESET_B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A4 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_Y (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1_N (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_Y (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A3 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A4 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_SET_B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_Y (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_B1_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap127_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SCD (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A1 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A4 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A4 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SCD (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A4 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_RESET_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A4 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_Y (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_B1_N (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SCD (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SET_B (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_B1_N (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_Y (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_B1_N (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_B1_N (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_Y (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_B1_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_Y (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_B1_N (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_Y (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SCE (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_Y (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_Y (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_D (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_S1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A3 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A3 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_Y (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1_N (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_Y (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SCE (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_Y (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_B1_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A3 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_X (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_D (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SCE (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A4 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_D (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_SET_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_B1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_Q (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_Q (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCE (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_Q (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_B1_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_X (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A4 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A4 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_X (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_SCD (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_X (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_Y (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A3 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SCE (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_X (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_D (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_Q (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_Q_N (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A3 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_Q (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_Y (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_S1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_B1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A3 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_Y (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_Y (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_D (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_X (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A3 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_S0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A0 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1_N (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCD (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_X (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A0 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A2 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_X (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A0 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_X (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_S0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A0 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A3 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A4 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_Q (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_X (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A4 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_SCE (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A3 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_X (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_X (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_S0 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCE (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SET_B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_SCE (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_Y (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1_N (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_Y (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCD (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_S0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_Y (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_S0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A3 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Y (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_X (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_B1_N (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A0 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_Y (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A0 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_B1 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_B1_N (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_X (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_X (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A0 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A3 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1_N (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B1_N (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A4 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_Y (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S0 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_D (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_X (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_S1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S0 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_X (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_RESET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_B1_N (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_X (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_X (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_X (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_s831_D (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_X (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_s842_D (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_X (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_X (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_X (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_RESET_B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A3 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_Y (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge782_A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge775_A3 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A0 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_B (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_Y (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_X (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_X (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S0 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_RESET_B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_X (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_Q (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_X (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_SCD (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_X (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_X (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B1_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCE (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_RESET_B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_B1_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire152_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_Y (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap150_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_Y (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_Q_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B1_N (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_Q (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_B1_N (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_B1_N (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_B (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_B1_N (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_Q (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_s809_Q (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_s811_Q (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A2 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_S1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A3 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net681_A (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_s812_GCLK (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_s818_Q (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S0 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_SET_B (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_s827_Q (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_B1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_B1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_Y (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_Q (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold50_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_Q (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_Y (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_Q (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_Q (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_S1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S0 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_Y (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_Y (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_SCD (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A4 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap135_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_D (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A4 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A4 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_Y (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_Y (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_Y (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_SCE (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_B1_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_A0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_Y (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A4 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Y (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_RESET_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_Y (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A4 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A4 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_SCE (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_B1_N (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCD (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S0 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A3 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_S0 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A4 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_SCD (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge766_SCE (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_B1_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_B1_N (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A0 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A4 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_D (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B1_N (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1_N (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_SCD (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A4 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_B1_N (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_B1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_RESET_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B1_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A0 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_A3 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A4 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SCD (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_SCE (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A2 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_B1_N (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_RESET_B (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_SCE (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_S0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_S0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_B1_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A3 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCD (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_B1_N (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A4 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A3 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A3 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_B1_N (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_SCD (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_B (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_B1_N (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_B1_N (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_B1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_B (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_D (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_SCE (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_B1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_B1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_S0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A0 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A4 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_B1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A4 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_S0 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A4 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A2 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_A3 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SCD (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A4 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B1_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_B1_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_SET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_B1_N (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B1_N (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A4 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_X (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_S1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge773_S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B1_N (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_X (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_B (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire130_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_B (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_Y (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_Y (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold46_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_B1_N (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A3 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S1 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A1 (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_Y (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_X (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S1 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_X (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_B1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_Y (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_SET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_B1_N (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A4 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_X (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S0 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_SCE (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_SET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_B1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_B1 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c124_B1_N (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_Y (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_Y (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A4 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_SCD (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_B1_N (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_SCD (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_SCE (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_B1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_Q (.DIODE(net875));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_X (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_SCD (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_B1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_X (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A4 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_SET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_B1 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_SET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A4 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_X (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_B1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_B1_N (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_SCE (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_B1 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B1_N (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S1 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A2 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_A4 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_SCE (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_SCE (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_SCE (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_SET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_A2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_SCE (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_B1_N (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_B1 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SCE (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B1_N (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_S0 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_RESET_B (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCE (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A4 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A4 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_SET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S0 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A3 (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_SCD (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B1_N (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A4 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A3 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_A4 (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_B1_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_B1_N (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap128_X (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_B1_N (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A4 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_B1_N (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_SCE (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire130_X (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_B1_N (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A4 (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_SET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A4 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_B1_N (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_B1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SCE (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap135_X (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_B1_N (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap136_X (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_A2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire137_X (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_B1 (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1_N (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A4 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A4 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_B1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_B1_N (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire141_X (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_B1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A2 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap144_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_B1_N (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_B1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap146_X (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_B1_N (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_B1 (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap149_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_D (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_B (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap150_X (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_X (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire152_X (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap151_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c111_B (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B1_N (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_S0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_SCD (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B1_N (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1_N (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1_N (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_B (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_SCD (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c85_B1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_B1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_A3 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_S1 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B1_N (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_B1_N (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_SET_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A4 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_X (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1_N (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s811_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s812_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_GATE_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s807_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_GATE (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s810_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s883_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s816_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s818_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s820_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s823_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s837_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge787_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s827_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s886_SLEEP_B (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s849_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s850_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s851_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s856_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s854_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s859_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s861_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s862_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s867_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s871_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s830_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s838_SLEEP_B (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s841_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s843_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s844_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s845_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s876_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s878_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S0 (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_B1 (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_S1 (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net682_X (.DIODE(clknet_1_0__leaf_net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S1 (.DIODE(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net681_X (.DIODE(clknet_1_0__leaf_net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_X (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_X (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer25_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer24_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer38_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer40_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer39_X (.DIODE(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer16 (.A(net93),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net211),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net987),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net837),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net989),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net990),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net837),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net992),
    .X(net993));
 sky130_fd_sc_hd__xnor2_1 clone47 (.A(net960),
    .B(net796),
    .Y(net994));
 sky130_fd_sc_hd__a21bo_1 clone48 (.A1(net827),
    .A2(net774),
    .B1_N(net773),
    .X(net995));
 sky130_fd_sc_hd__a21bo_1 clone49 (.A1(net909),
    .A2(net77),
    .B1_N(net635),
    .X(net996));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer50 (.A(net77),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net997),
    .X(net998));
 sky130_fd_sc_hd__a21bo_1 clone52 (.A1(net894),
    .A2(net194),
    .B1_N(net895),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net65),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net321),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net321),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net1002),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net321),
    .X(net1004));
 sky130_fd_sc_hd__a21bo_1 clone58 (.A1(net827),
    .A2(net774),
    .B1_N(net773),
    .X(net1005));
 sky130_fd_sc_hd__xnor2_1 clone59 (.A(net71),
    .B(net64),
    .Y(net1006));
 sky130_fd_sc_hd__clkbuf_1 clone60 (.A(net885),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_1 clone61 (.A(net63),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net118),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net118),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net118),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net118),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net118),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(net1013),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(net201),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(net1015),
    .X(net1016));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer70 (.A(net1016),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net1017),
    .X(net1018));
 sky130_fd_sc_hd__xnor2_1 clone72 (.A(net96),
    .B(net210),
    .Y(net1019));
 sky130_fd_sc_hd__clkbuf_1 clone73 (.A(net76),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_1 clone74 (.A(net61),
    .X(net1021));
 sky130_fd_sc_hd__xnor2_1 clone75 (.A(net70),
    .B(net812),
    .Y(net1022));
 sky130_fd_sc_hd__clkbuf_1 clone76 (.A(net333),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net812),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net885),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer79 (.A(net1025),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net1025),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer81 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer82 (.A(net92),
    .X(net1029));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
