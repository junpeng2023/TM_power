module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in62,
    in63,
    in64,
    in65,
    in66,
    in67,
    in68,
    in69,
    in7,
    in70,
    in71,
    in72,
    in73,
    in74,
    in75,
    in76,
    in77,
    in78,
    in79,
    in8,
    in80,
    in81,
    in82,
    in83,
    in84,
    in85,
    in86,
    in87,
    in88,
    in89,
    in9,
    in90,
    in91,
    in92,
    in93,
    in94,
    in95,
    in96,
    in97,
    in98,
    in99,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out62,
    out63,
    out64,
    out65,
    out66,
    out67,
    out68,
    out69,
    out7,
    out70,
    out71,
    out72,
    out73,
    out74,
    out75,
    out76,
    out77,
    out78,
    out79,
    out8,
    out80,
    out81,
    out82,
    out83,
    out84,
    out85,
    out86,
    out87,
    out88,
    out89,
    out9,
    out90,
    out91,
    out92,
    out93,
    out94,
    out95,
    out96,
    out97,
    out98,
    out99,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in62;
 input in63;
 input in64;
 input in65;
 input in66;
 input in67;
 input in68;
 input in69;
 input in7;
 input in70;
 input in71;
 input in72;
 input in73;
 input in74;
 input in75;
 input in76;
 input in77;
 input in78;
 input in79;
 input in8;
 input in80;
 input in81;
 input in82;
 input in83;
 input in84;
 input in85;
 input in86;
 input in87;
 input in88;
 input in89;
 input in9;
 input in90;
 input in91;
 input in92;
 input in93;
 input in94;
 input in95;
 input in96;
 input in97;
 input in98;
 input in99;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out62;
 output out63;
 output out64;
 output out65;
 output out66;
 output out67;
 output out68;
 output out69;
 output out7;
 output out70;
 output out71;
 output out72;
 output out73;
 output out74;
 output out75;
 output out76;
 output out77;
 output out78;
 output out79;
 output out8;
 output out80;
 output out81;
 output out82;
 output out83;
 output out84;
 output out85;
 output out86;
 output out87;
 output out88;
 output out89;
 output out9;
 output out90;
 output out91;
 output out92;
 output out93;
 output out94;
 output out95;
 output out96;
 output out97;
 output out98;
 output out99;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net39;
 wire net167;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net754;
 wire clknet_1_0__leaf_net754;
 wire clknet_1_1__leaf_net754;
 wire clknet_0_net467;
 wire clknet_1_0__leaf_net467;
 wire clknet_1_1__leaf_net467;
 wire clknet_0_net753;
 wire clknet_1_0__leaf_net753;
 wire clknet_1_1__leaf_net753;
 wire clknet_0_net752;
 wire clknet_1_0__leaf_net752;
 wire clknet_1_1__leaf_net752;
 wire clknet_0_net734;
 wire clknet_1_0__leaf_net734;
 wire clknet_1_1__leaf_net734;
 wire clknet_0_net733;
 wire clknet_1_0__leaf_net733;
 wire clknet_1_1__leaf_net733;
 wire clknet_0_net732;
 wire clknet_1_0__leaf_net732;
 wire clknet_1_1__leaf_net732;
 wire clknet_0_net452;
 wire clknet_1_0__leaf_net452;
 wire clknet_1_1__leaf_net452;
 wire clknet_0_net476;
 wire clknet_1_0__leaf_net476;
 wire clknet_1_1__leaf_net476;
 wire clknet_0_net446;
 wire clknet_1_0__leaf_net446;
 wire clknet_1_1__leaf_net446;
 wire clknet_0_net696;
 wire clknet_1_0__leaf_net696;
 wire clknet_1_1__leaf_net696;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net676;
 wire clknet_1_0__leaf_net676;
 wire clknet_1_1__leaf_net676;
 wire clknet_0_net417;
 wire clknet_1_0__leaf_net417;
 wire clknet_1_1__leaf_net417;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net416;
 wire clknet_1_0__leaf_net416;
 wire clknet_1_1__leaf_net416;
 wire clknet_0_net346;
 wire clknet_1_0__leaf_net346;
 wire clknet_1_1__leaf_net346;
 wire clknet_0_net349;
 wire clknet_1_0__leaf_net349;
 wire clknet_1_1__leaf_net349;
 wire clknet_0_net339;
 wire clknet_1_0__leaf_net339;
 wire clknet_1_1__leaf_net339;
 wire clknet_0_net348;
 wire clknet_1_0__leaf_net348;
 wire clknet_1_1__leaf_net348;
 wire clknet_0_net888;
 wire clknet_1_0__leaf_net888;
 wire clknet_1_1__leaf_net888;
 wire clknet_0_net444;
 wire clknet_1_0__leaf_net444;
 wire clknet_1_1__leaf_net444;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net428;
 wire clknet_1_0__leaf_net428;
 wire clknet_1_1__leaf_net428;
 wire clknet_0_net418;
 wire clknet_1_0__leaf_net418;
 wire clknet_1_1__leaf_net418;
 wire clknet_0_net367;
 wire clknet_1_0__leaf_net367;
 wire clknet_1_1__leaf_net367;
 wire clknet_0_net372;
 wire clknet_1_0__leaf_net372;
 wire clknet_1_1__leaf_net372;
 wire clknet_0_net675;
 wire clknet_1_0__leaf_net675;
 wire clknet_1_1__leaf_net675;
 wire clknet_0_net324;
 wire clknet_1_0__leaf_net324;
 wire clknet_1_1__leaf_net324;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net638;
 wire clknet_1_0__leaf_net638;
 wire clknet_1_1__leaf_net638;
 wire clknet_0_net357;
 wire clknet_1_0__leaf_net357;
 wire clknet_1_1__leaf_net357;
 wire clknet_0_net637;
 wire clknet_1_0__leaf_net637;
 wire clknet_1_1__leaf_net637;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net261;
 wire clknet_1_0__leaf_net261;
 wire clknet_1_1__leaf_net261;
 wire clknet_0_net258;
 wire clknet_1_0__leaf_net258;
 wire clknet_1_1__leaf_net258;
 wire clknet_0_net257;
 wire clknet_1_0__leaf_net257;
 wire clknet_1_1__leaf_net257;
 wire clknet_0_net890;
 wire clknet_1_0__leaf_net890;
 wire clknet_1_1__leaf_net890;
 wire clknet_0_net618;
 wire clknet_1_0__leaf_net618;
 wire clknet_1_1__leaf_net618;
 wire clknet_0_net388;
 wire clknet_1_0__leaf_net388;
 wire clknet_1_1__leaf_net388;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net617;
 wire clknet_1_0__leaf_net617;
 wire clknet_1_1__leaf_net617;
 wire clknet_0_net313;
 wire clknet_1_0__leaf_net313;
 wire clknet_1_1__leaf_net313;
 wire clknet_0_net616;
 wire clknet_1_0__leaf_net616;
 wire clknet_1_1__leaf_net616;
 wire clknet_0_net598;
 wire clknet_1_0__leaf_net598;
 wire clknet_1_1__leaf_net598;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net241;
 wire clknet_1_0__leaf_net241;
 wire clknet_1_1__leaf_net241;
 wire clknet_0_net240;
 wire clknet_1_0__leaf_net240;
 wire clknet_1_1__leaf_net240;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net329;
 wire clknet_1_0__leaf_net329;
 wire clknet_1_1__leaf_net329;
 wire clknet_0_net204;
 wire clknet_1_0__leaf_net204;
 wire clknet_1_1__leaf_net204;
 wire clknet_0_net411;
 wire clknet_1_0__leaf_net411;
 wire clknet_1_1__leaf_net411;
 wire clknet_0_net399;
 wire clknet_1_0__leaf_net399;
 wire clknet_1_1__leaf_net399;
 wire clknet_0_net340;
 wire clknet_1_0__leaf_net340;
 wire clknet_1_1__leaf_net340;
 wire clknet_0_net312;
 wire clknet_1_0__leaf_net312;
 wire clknet_1_1__leaf_net312;
 wire clknet_0_net581;
 wire clknet_1_0__leaf_net581;
 wire clknet_1_1__leaf_net581;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net580;
 wire clknet_1_0__leaf_net580;
 wire clknet_1_1__leaf_net580;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net918;
 wire clknet_1_0__leaf_net918;
 wire clknet_1_1__leaf_net918;
 wire clknet_0_net563;
 wire clknet_1_0__leaf_net563;
 wire clknet_1_1__leaf_net563;
 wire clknet_0_net247;
 wire clknet_1_0__leaf_net247;
 wire clknet_1_1__leaf_net247;
 wire clknet_0_net148;
 wire clknet_1_0__leaf_net148;
 wire clknet_1_1__leaf_net148;
 wire clknet_0_net884;
 wire clknet_1_0__leaf_net884;
 wire clknet_1_1__leaf_net884;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net229;
 wire clknet_1_0__leaf_net229;
 wire clknet_1_1__leaf_net229;
 wire clknet_0_net337;
 wire clknet_1_0__leaf_net337;
 wire clknet_1_1__leaf_net337;
 wire clknet_0_net342;
 wire clknet_1_0__leaf_net342;
 wire clknet_1_1__leaf_net342;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net893;
 wire clknet_1_0__leaf_net893;
 wire clknet_1_1__leaf_net893;
 wire clknet_0_net280;
 wire clknet_1_0__leaf_net280;
 wire clknet_1_1__leaf_net280;
 wire clknet_0_net282;
 wire clknet_1_0__leaf_net282;
 wire clknet_1_1__leaf_net282;
 wire clknet_0_net141;
 wire clknet_1_0__leaf_net141;
 wire clknet_1_1__leaf_net141;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net147;
 wire clknet_1_0__leaf_net147;
 wire clknet_1_1__leaf_net147;
 wire clknet_0_net156;
 wire clknet_1_0__leaf_net156;
 wire clknet_1_1__leaf_net156;
 wire clknet_0_net159;
 wire clknet_1_0__leaf_net159;
 wire clknet_1_1__leaf_net159;
 wire clknet_0_net908;
 wire clknet_1_0__leaf_net908;
 wire clknet_1_1__leaf_net908;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net870;
 wire clknet_1_0__leaf_net870;
 wire clknet_1_1__leaf_net870;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net136;
 wire clknet_1_0__leaf_net136;
 wire clknet_1_1__leaf_net136;
 wire clknet_0_net544;
 wire clknet_1_0__leaf_net544;
 wire clknet_1_1__leaf_net544;
 wire clknet_0_net363;
 wire clknet_1_0__leaf_net363;
 wire clknet_1_1__leaf_net363;
 wire clknet_0_net291;
 wire clknet_1_0__leaf_net291;
 wire clknet_1_1__leaf_net291;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net405;
 wire clknet_1_0__leaf_net405;
 wire clknet_1_1__leaf_net405;
 wire clknet_0_net397;
 wire clknet_1_0__leaf_net397;
 wire clknet_1_1__leaf_net397;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net415;
 wire clknet_1_0__leaf_net415;
 wire clknet_1_1__leaf_net415;
 wire clknet_0_net409;
 wire clknet_1_0__leaf_net409;
 wire clknet_1_1__leaf_net409;
 wire clknet_0_net396;
 wire clknet_1_0__leaf_net396;
 wire clknet_1_1__leaf_net396;
 wire clknet_0_net408;
 wire clknet_1_0__leaf_net408;
 wire clknet_1_1__leaf_net408;
 wire clknet_0_net297;
 wire clknet_1_0__leaf_net297;
 wire clknet_1_1__leaf_net297;
 wire clknet_0_net299;
 wire clknet_1_0__leaf_net299;
 wire clknet_1_1__leaf_net299;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net295;
 wire clknet_1_0__leaf_net295;
 wire clknet_1_1__leaf_net295;
 wire clknet_0_net131;
 wire clknet_1_0__leaf_net131;
 wire clknet_1_1__leaf_net131;
 wire clknet_0_net132;
 wire clknet_1_0__leaf_net132;
 wire clknet_1_1__leaf_net132;
 wire clknet_0_net883;
 wire clknet_1_0__leaf_net883;
 wire clknet_1_1__leaf_net883;
 wire clknet_0_net112;
 wire clknet_1_0__leaf_net112;
 wire clknet_1_1__leaf_net112;
 wire clknet_0_net114;
 wire clknet_1_0__leaf_net114;
 wire clknet_1_1__leaf_net114;
 wire clknet_0_net133;
 wire clknet_1_0__leaf_net133;
 wire clknet_1_1__leaf_net133;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net899;
 wire clknet_1_0__leaf_net899;
 wire clknet_1_1__leaf_net899;
 wire clknet_0_net116;
 wire clknet_1_0__leaf_net116;
 wire clknet_1_1__leaf_net116;
 wire clknet_0_net122;
 wire clknet_1_0__leaf_net122;
 wire clknet_1_1__leaf_net122;
 wire clknet_0_net115;
 wire clknet_1_0__leaf_net115;
 wire clknet_1_1__leaf_net115;
 wire clknet_0_net278;
 wire clknet_1_0__leaf_net278;
 wire clknet_1_1__leaf_net278;
 wire clknet_0_net543;
 wire clknet_1_0__leaf_net543;
 wire clknet_1_1__leaf_net543;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net207;
 wire clknet_1_0__leaf_net207;
 wire clknet_1_1__leaf_net207;
 wire clknet_0_net429;
 wire clknet_1_0__leaf_net429;
 wire clknet_1_1__leaf_net429;
 wire clknet_0_net220;
 wire clknet_1_0__leaf_net220;
 wire clknet_1_1__leaf_net220;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net194;
 wire clknet_1_0__leaf_net194;
 wire clknet_1_1__leaf_net194;
 wire clknet_0_net111;
 wire clknet_1_0__leaf_net111;
 wire clknet_1_1__leaf_net111;
 wire clknet_0_net542;
 wire clknet_1_0__leaf_net542;
 wire clknet_1_1__leaf_net542;
 wire clknet_0_net529;
 wire clknet_1_0__leaf_net529;
 wire clknet_1_1__leaf_net529;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net904;
 wire clknet_1_0__leaf_net904;
 wire clknet_1_1__leaf_net904;
 wire clknet_0_net885;
 wire clknet_1_0__leaf_net885;
 wire clknet_1_1__leaf_net885;
 wire clknet_0_net83;
 wire clknet_1_0__leaf_net83;
 wire clknet_1_1__leaf_net83;
 wire clknet_0_net56;
 wire clknet_1_0__leaf_net56;
 wire clknet_1_1__leaf_net56;
 wire clknet_0_net62;
 wire clknet_1_0__leaf_net62;
 wire clknet_1_1__leaf_net62;
 wire clknet_0_net59;
 wire clknet_1_0__leaf_net59;
 wire clknet_1_1__leaf_net59;
 wire clknet_0_net254;
 wire clknet_1_0__leaf_net254;
 wire clknet_1_1__leaf_net254;
 wire clknet_0_net253;
 wire clknet_1_0__leaf_net253;
 wire clknet_1_1__leaf_net253;
 wire clknet_0_net248;
 wire clknet_1_0__leaf_net248;
 wire clknet_1_1__leaf_net248;
 wire clknet_0_net920;
 wire clknet_1_0__leaf_net920;
 wire clknet_1_1__leaf_net920;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net927;
 wire clknet_1_0__leaf_net927;
 wire clknet_1_1__leaf_net927;
 wire clknet_0_net64;
 wire clknet_1_0__leaf_net64;
 wire clknet_1_1__leaf_net64;
 wire clknet_0_net61;
 wire clknet_1_0__leaf_net61;
 wire clknet_1_1__leaf_net61;
 wire clknet_0_net57;
 wire clknet_1_0__leaf_net57;
 wire clknet_1_1__leaf_net57;
 wire clknet_0_net78;
 wire clknet_1_0__leaf_net78;
 wire clknet_1_1__leaf_net78;
 wire clknet_0_net923;
 wire clknet_1_0__leaf_net923;
 wire clknet_1_1__leaf_net923;
 wire clknet_0_net75;
 wire clknet_1_0__leaf_net75;
 wire clknet_1_1__leaf_net75;
 wire clknet_0_net916;
 wire clknet_1_0__leaf_net916;
 wire clknet_1_1__leaf_net916;
 wire clknet_0_net528;
 wire clknet_1_0__leaf_net528;
 wire clknet_1_1__leaf_net528;
 wire clknet_0_net158;
 wire clknet_1_0__leaf_net158;
 wire clknet_1_1__leaf_net158;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net160;
 wire clknet_1_0__leaf_net160;
 wire clknet_1_1__leaf_net160;
 wire clknet_0_net47;
 wire clknet_1_0__leaf_net47;
 wire clknet_1_1__leaf_net47;
 wire clknet_0_net882;
 wire clknet_1_0__leaf_net882;
 wire clknet_1_1__leaf_net882;
 wire clknet_0_net243;
 wire clknet_1_0__leaf_net243;
 wire clknet_1_1__leaf_net243;
 wire clknet_0_net73;
 wire clknet_1_0__leaf_net73;
 wire clknet_1_1__leaf_net73;
 wire clknet_0_net54;
 wire clknet_1_0__leaf_net54;
 wire clknet_1_1__leaf_net54;
 wire clknet_0_net137;
 wire clknet_1_0__leaf_net137;
 wire clknet_1_1__leaf_net137;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;

 sky130_fd_sc_hd__mux4_1 c100 (.A0(net856),
    .A1(net868),
    .A2(net852),
    .A3(net865),
    .S0(net851),
    .S1(net853),
    .X(net0));
 sky130_fd_sc_hd__mux4_2 c101 (.A0(net792),
    .A1(net788),
    .A2(net786),
    .A3(net867),
    .S0(net807),
    .S1(net868),
    .X(net910));
 sky130_fd_sc_hd__mux4_2 c102 (.A0(net786),
    .A1(net1010),
    .A2(net790),
    .A3(net1011),
    .S0(net868),
    .S1(net852),
    .X(net1));
 sky130_fd_sc_hd__mux4_2 c103 (.A0(net852),
    .A1(net986),
    .A2(net1),
    .A3(net853),
    .S0(net837),
    .S1(net829),
    .X(net2));
 sky130_fd_sc_hd__mux4_2 c104 (.A0(net860),
    .A1(net2),
    .A2(net855),
    .A3(net842),
    .S0(net1),
    .S1(net820),
    .X(net939));
 sky130_fd_sc_hd__mux4_2 c116 (.A0(net829),
    .A1(net855),
    .A2(net939),
    .A3(net800),
    .S0(net1010),
    .S1(net857),
    .X(net940));
 sky130_fd_sc_hd__mux4_1 c117 (.A0(net1002),
    .A1(net796),
    .A2(net940),
    .A3(net829),
    .S0(net810),
    .S1(net863),
    .X(net3));
 sky130_fd_sc_hd__mux4_2 c118 (.A0(net3),
    .A1(net1011),
    .A2(net843),
    .A3(net850),
    .S0(net997),
    .S1(net796),
    .X(net924));
 sky130_fd_sc_hd__mux4_2 c119 (.A0(net842),
    .A1(net804),
    .A2(net867),
    .A3(net834),
    .S0(net850),
    .S1(net924),
    .X(net936));
 sky130_fd_sc_hd__mux4_2 c120 (.A0(net850),
    .A1(net940),
    .A2(net792),
    .A3(net924),
    .S0(net867),
    .S1(net939),
    .X(net934));
 sky130_fd_sc_hd__mux4_2 c121 (.A0(net796),
    .A1(net3),
    .A2(net934),
    .A3(net924),
    .S0(net863),
    .S1(net862),
    .X(net922));
 sky130_fd_sc_hd__mux4_2 c122 (.A0(net863),
    .A1(net924),
    .A2(net934),
    .A3(net850),
    .S0(net922),
    .S1(net936),
    .X(net937));
 sky130_fd_sc_hd__mux4_2 c123 (.A0(net778),
    .A1(net937),
    .A2(net855),
    .A3(net924),
    .S0(net922),
    .S1(net934),
    .X(net938));
 sky130_fd_sc_hd__mux4_1 c124 (.A0(net3),
    .A1(net936),
    .A2(net938),
    .A3(net829),
    .S0(net940),
    .S1(net922),
    .X(net896));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net800),
    .A1(net938),
    .A2(net896),
    .A3(net937),
    .S0(net867),
    .S1(net924),
    .X(net935));
 sky130_fd_sc_hd__a41o_4 c126 (.A1(net1074),
    .A2(net814),
    .A3(net167),
    .A4(net990),
    .B1(net996),
    .X(net4));
 sky130_fd_sc_hd__mux4_2 c127 (.A0(net999),
    .A1(net983),
    .A2(net994),
    .A3(net990),
    .S0(net996),
    .S1(net1071),
    .X(net5));
 sky130_fd_sc_hd__a41o_4 c128 (.A1(net5),
    .A2(net792),
    .A3(net778),
    .A4(net1002),
    .B1(net983),
    .X(net921));
 sky130_fd_sc_hd__a41o_4 c129 (.A1(net978),
    .A2(net990),
    .A3(net979),
    .A4(net983),
    .B1(net1002),
    .X(net6));
 sky130_fd_sc_hd__a41o_4 c130 (.A1(net1072),
    .A2(net1018),
    .A3(net978),
    .A4(net983),
    .B1(net976),
    .X(net7));
 sky130_fd_sc_hd__a41o_4 c131 (.A1(net975),
    .A2(net978),
    .A3(net979),
    .A4(net1002),
    .B1(net996),
    .X(net8));
 sky130_fd_sc_hd__a41o_4 c132 (.A1(net974),
    .A2(net1075),
    .A3(net979),
    .A4(net990),
    .B1(net975),
    .X(net9));
 sky130_fd_sc_hd__mux4_2 c133 (.A0(net976),
    .A1(net979),
    .A2(net970),
    .A3(net1008),
    .S0(net975),
    .S1(net792),
    .X(net10));
 sky130_fd_sc_hd__mux4_2 c134 (.A0(net167),
    .A1(net778),
    .A2(net974),
    .A3(net979),
    .S0(net970),
    .S1(net966),
    .X(net11));
 sky130_fd_sc_hd__mux4_2 c135 (.A0(net976),
    .A1(net975),
    .A2(net1015),
    .A3(net978),
    .S0(net965),
    .S1(net967),
    .X(net12));
 sky130_fd_sc_hd__mux4_2 c136 (.A0(net976),
    .A1(net964),
    .A2(net996),
    .A3(net965),
    .S0(net974),
    .S1(net1071),
    .X(net13));
 sky130_fd_sc_hd__mux4_2 c137 (.A0(net13),
    .A1(net965),
    .A2(net778),
    .A3(net1011),
    .S0(net1059),
    .S1(net970),
    .X(net14));
 sky130_fd_sc_hd__mux4_2 c138 (.A0(net1071),
    .A1(net13),
    .A2(net966),
    .A3(net1072),
    .S0(net996),
    .S1(net974),
    .X(net15));
 sky130_fd_sc_hd__mux4_2 c139 (.A0(net15),
    .A1(net990),
    .A2(net792),
    .A3(net167),
    .S0(net966),
    .S1(net13),
    .X(net16));
 sky130_fd_sc_hd__mux4_2 c140 (.A0(net958),
    .A1(net15),
    .A2(net1000),
    .A3(net990),
    .S0(net976),
    .S1(net978),
    .X(net17));
 sky130_fd_sc_hd__mux4_2 c141 (.A0(net1049),
    .A1(net17),
    .A2(net15),
    .A3(net13),
    .S0(net958),
    .S1(net966),
    .X(net18));
 sky130_fd_sc_hd__mux4_2 c142 (.A0(net1074),
    .A1(net17),
    .A2(net15),
    .A3(net1072),
    .S0(net18),
    .S1(net958),
    .X(net19));
 sky130_fd_sc_hd__mux4_2 c143 (.A0(net17),
    .A1(net964),
    .A2(net15),
    .A3(net970),
    .S0(net958),
    .S1(net1024),
    .X(net926));
 sky130_fd_sc_hd__mux4_2 c144 (.A0(net970),
    .A1(net17),
    .A2(net19),
    .A3(net1024),
    .S0(net926),
    .S1(net18),
    .X(net915));
 sky130_fd_sc_hd__mux4_2 c145 (.A0(net1059),
    .A1(net926),
    .A2(net1084),
    .A3(net949),
    .S0(net964),
    .S1(net1055),
    .X(net20));
 sky130_fd_sc_hd__mux4_2 c146 (.A0(net1024),
    .A1(net1050),
    .A2(net20),
    .A3(net1084),
    .S0(net1021),
    .S1(net926),
    .X(net21));
 sky130_fd_sc_hd__a41o_1 c147 (.A1(net1018),
    .A2(net979),
    .A3(net921),
    .A4(net975),
    .B1(net788),
    .X(net22));
 sky130_fd_sc_hd__mux4_2 c148 (.A0(net792),
    .A1(net789),
    .A2(net1009),
    .A3(net17),
    .S0(net1069),
    .S1(net784),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 c149 (.A0(net1069),
    .A1(net793),
    .A2(net789),
    .A3(net990),
    .S0(net1011),
    .S1(net794),
    .X(net912));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net794),
    .A1(net814),
    .A2(net793),
    .A3(net1067),
    .S0(net921),
    .S1(net23),
    .X(net24));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net804),
    .A1(net1069),
    .A2(net1074),
    .A3(net789),
    .S0(net1073),
    .S1(net950),
    .X(net25));
 sky130_fd_sc_hd__mux4_2 c152 (.A0(net784),
    .A1(net795),
    .A2(net9),
    .A3(net799),
    .S0(net1072),
    .S1(net1069),
    .X(net932));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net1009),
    .A1(net5),
    .A2(net792),
    .A3(net814),
    .S0(net789),
    .S1(net794),
    .X(net26));
 sky130_fd_sc_hd__mux4_2 c154 (.A0(net1067),
    .A1(net25),
    .A2(net966),
    .A3(net1068),
    .S0(net1070),
    .S1(net1075),
    .X(net27));
 sky130_fd_sc_hd__mux4_2 c155 (.A0(net1070),
    .A1(net794),
    .A2(net13),
    .A3(net27),
    .S0(net25),
    .S1(net1069),
    .X(net28));
 sky130_fd_sc_hd__mux4_2 c156 (.A0(net795),
    .A1(net950),
    .A2(net28),
    .A3(net1070),
    .S0(net23),
    .S1(net27),
    .X(net29));
 sky130_fd_sc_hd__mux4_2 c157 (.A0(net27),
    .A1(net795),
    .A2(net25),
    .A3(net948),
    .S0(net1069),
    .S1(net994),
    .X(net894));
 sky130_fd_sc_hd__mux4_1 c158 (.A0(net1026),
    .A1(net1068),
    .A2(net1002),
    .A3(net1035),
    .S0(net1023),
    .S1(net1071),
    .X(net30));
 sky130_fd_sc_hd__mux4_2 c159 (.A0(net794),
    .A1(net814),
    .A2(net28),
    .A3(net25),
    .S0(net1070),
    .S1(net1069),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 c160 (.A0(net31),
    .A1(net1020),
    .A2(net1010),
    .A3(net1067),
    .S0(net1035),
    .S1(net1059),
    .X(net32));
 sky130_fd_sc_hd__mux4_2 c161 (.A0(net31),
    .A1(net1070),
    .A2(net926),
    .A3(net19),
    .S0(net950),
    .S1(net524),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 c162 (.A0(net1050),
    .A1(net1026),
    .A2(net33),
    .A3(net1009),
    .S0(net1046),
    .S1(net523),
    .X(net34));
 sky130_fd_sc_hd__mux4_1 c163 (.A0(net1022),
    .A1(net1032),
    .A2(net778),
    .A3(net33),
    .S0(net522),
    .S1(net525),
    .X(net35));
 sky130_fd_sc_hd__mux4_2 c164 (.A0(net1008),
    .A1(net1020),
    .A2(net20),
    .A3(net1067),
    .S0(net525),
    .S1(net526),
    .X(net36));
 sky130_fd_sc_hd__mux4_2 c165 (.A0(net1046),
    .A1(net1022),
    .A2(net31),
    .A3(net1068),
    .S0(net948),
    .S1(net526),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c166 (.A0(net946),
    .A1(net943),
    .A2(net1068),
    .A3(net1041),
    .S0(net33),
    .S1(net1063),
    .X(net38));
 sky130_fd_sc_hd__mux4_2 c167 (.A0(net1068),
    .A1(net33),
    .A2(net799),
    .A3(net944),
    .S1(net526),
    .X(net513));
 sky130_fd_sc_hd__mux4_2 c168 (.A0(net823),
    .A1(net23),
    .A2(net800),
    .A3(net1068),
    .S0(net811),
    .S1(net1072),
    .X(net40));
 sky130_fd_sc_hd__mux4_2 c169 (.A0(net806),
    .A1(net822),
    .A2(net40),
    .A3(net1041),
    .S0(net823),
    .S1(net946),
    .X(net41));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net979),
    .A1(net817),
    .A2(net791),
    .A3(net1073),
    .S0(net821),
    .S1(net804),
    .X(net42));
 sky130_fd_sc_hd__mux4_2 c171 (.A0(net1074),
    .A1(net784),
    .A2(net42),
    .A3(net1010),
    .S0(net808),
    .S1(net991),
    .X(net43));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(net41),
    .A1(net1046),
    .A2(net18),
    .A3(net783),
    .S0(net43),
    .S1(net819),
    .X(net44));
 sky130_fd_sc_hd__mux4_1 c173 (.A0(net41),
    .A1(net788),
    .A2(net1023),
    .A3(net797),
    .S0(net822),
    .S1(net527),
    .X(net45));
 sky130_fd_sc_hd__mux4_2 c174 (.A0(net811),
    .A1(net42),
    .A2(net40),
    .A3(net817),
    .S0(net804),
    .S1(net526),
    .X(net46));
 sky130_fd_sc_hd__mux4_1 c175 (.A0(net42),
    .A1(net1003),
    .A2(net1009),
    .A3(net1073),
    .S0(net818),
    .S1(clknet_1_1__leaf_net528),
    .X(net47));
 sky130_fd_sc_hd__mux4_2 c176 (.A0(net783),
    .A1(net819),
    .A2(net817),
    .A3(net984),
    .S0(net926),
    .S1(net1067),
    .X(net48));
 sky130_fd_sc_hd__mux4_2 c177 (.A0(net824),
    .A1(net807),
    .A2(net806),
    .A3(net962),
    .S0(net522),
    .S1(net527),
    .X(net49));
 sky130_fd_sc_hd__mux4_2 c178 (.A0(net962),
    .A1(net18),
    .A2(net812),
    .A3(net1071),
    .S0(net20),
    .S1(net946),
    .X(net50));
 sky130_fd_sc_hd__mux4_1 c179 (.A0(net778),
    .A1(net50),
    .A2(net826),
    .A3(net41),
    .S0(net40),
    .S1(clknet_1_1__leaf_net528),
    .X(net51));
 sky130_fd_sc_hd__mux4_2 c180 (.A0(net819),
    .A1(net811),
    .A2(net1003),
    .A3(net48),
    .S0(net49),
    .S1(net806),
    .X(net52));
 sky130_fd_sc_hd__mux4_1 c181 (.A0(net18),
    .A1(net818),
    .A2(net49),
    .A3(net946),
    .S0(clknet_1_0__leaf_net47),
    .S1(clknet_1_0__leaf_net898),
    .X(net916));
 sky130_fd_sc_hd__mux4_1 c182 (.A0(net1084),
    .A1(net1006),
    .A2(net42),
    .A3(net48),
    .S0(net800),
    .S1(clknet_1_0__leaf_net47),
    .X(net882));
 sky130_fd_sc_hd__mux4_1 c183 (.A0(net812),
    .A1(net42),
    .A2(net43),
    .A3(net50),
    .S0(net784),
    .S1(clknet_1_1__leaf_net528),
    .X(net53));
 sky130_fd_sc_hd__mux4_1 c184 (.A0(net43),
    .A1(net1009),
    .A2(net793),
    .A3(clknet_1_1__leaf_net882),
    .S0(net1069),
    .S1(net1049),
    .X(net54));
 sky130_fd_sc_hd__mux4_1 c185 (.A0(net49),
    .A1(net949),
    .A2(net991),
    .A3(clknet_1_0__leaf_net54),
    .S0(clknet_1_1__leaf_net916),
    .S1(net527),
    .X(net55));
 sky130_fd_sc_hd__mux4_1 c186 (.A0(clknet_1_0__leaf_net47),
    .A1(net48),
    .A2(net46),
    .A3(net40),
    .S0(net43),
    .S1(clknet_1_0__leaf_net898),
    .X(net56));
 sky130_fd_sc_hd__mux4_1 c187 (.A0(clknet_1_1__leaf_net56),
    .A1(net812),
    .A2(net799),
    .A3(net811),
    .S0(net19),
    .S1(net508),
    .X(net57));
 sky130_fd_sc_hd__mux4_1 c188 (.A0(clknet_1_1__leaf_net916),
    .A1(clknet_1_1__leaf_net882),
    .A2(net20),
    .A3(net788),
    .S0(clknet_1_1__leaf_net57),
    .S1(net507),
    .X(net58));
 sky130_fd_sc_hd__mux4_2 c189 (.A0(net20),
    .A1(net1003),
    .A2(net1010),
    .A3(net967),
    .S0(clknet_1_1__leaf_net56),
    .S1(net513),
    .X(net59));
 sky130_fd_sc_hd__mux4_1 c190 (.A0(clknet_1_1__leaf_net59),
    .A1(net1073),
    .A2(net816),
    .A3(net20),
    .S0(clknet_1_0__leaf_net916),
    .S1(net946),
    .X(net60));
 sky130_fd_sc_hd__mux4_2 c191 (.A0(net1025),
    .A1(net837),
    .A2(net1019),
    .A3(net823),
    .S0(net845),
    .S1(net1009),
    .X(net906));
 sky130_fd_sc_hd__mux4_2 c192 (.A0(net42),
    .A1(net834),
    .A2(net1068),
    .A3(clknet_1_0__leaf_net59),
    .S0(net818),
    .S1(net48),
    .X(net61));
 sky130_fd_sc_hd__mux4_1 c193 (.A0(net49),
    .A1(net839),
    .A2(net25),
    .A3(net1061),
    .S0(net23),
    .S1(net517),
    .X(net927));
 sky130_fd_sc_hd__mux4_2 c194 (.A0(clknet_1_0__leaf_net56),
    .A1(clknet_1_0__leaf_net47),
    .A2(net986),
    .A3(net838),
    .S0(clknet_1_1__leaf_net61),
    .S1(net1062),
    .X(net62));
 sky130_fd_sc_hd__mux4_1 c195 (.A0(net832),
    .A1(net1032),
    .A2(clknet_1_1__leaf_net61),
    .A3(clknet_1_0__leaf_net56),
    .S0(net835),
    .S1(net50),
    .X(net63));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(clknet_1_1__leaf_net927),
    .A1(net820),
    .A2(net986),
    .A3(net849),
    .S0(net819),
    .S1(net1051),
    .X(net64));
 sky130_fd_sc_hd__mux4_1 c197 (.A0(net20),
    .A1(clknet_1_0__leaf_net61),
    .A2(net795),
    .A3(net1073),
    .S0(clknet_1_0__leaf_net59),
    .S1(net1003),
    .X(net931));
 sky130_fd_sc_hd__mux4_1 c198 (.A0(net824),
    .A1(net21),
    .A2(clknet_1_1__leaf_net61),
    .A3(net846),
    .S0(net1061),
    .S1(clknet_1_0__leaf_net62),
    .X(net65));
 sky130_fd_sc_hd__mux4_1 c199 (.A0(net943),
    .A1(net824),
    .A2(net21),
    .A3(clknet_1_1__leaf_net528),
    .S0(net933),
    .S1(net531),
    .X(net66));
 sky130_fd_sc_hd__mux4_2 c200 (.A0(net23),
    .A1(net1006),
    .A2(net787),
    .A3(net513),
    .S0(net530),
    .S1(net531),
    .X(net67));
 sky130_fd_sc_hd__mux4_1 c201 (.A0(clknet_1_1__leaf_net931),
    .A1(net792),
    .A2(net835),
    .A3(net941),
    .S0(net1009),
    .S1(net532),
    .X(net68));
 sky130_fd_sc_hd__mux4_1 c202 (.A0(clknet_1_0__leaf_net59),
    .A1(net906),
    .A2(net1068),
    .A3(clknet_1_0__leaf_net61),
    .S0(net832),
    .S1(net534),
    .X(net920));
 sky130_fd_sc_hd__mux4_1 c203 (.A0(net999),
    .A1(clknet_1_1__leaf_net920),
    .A2(clknet_1_0__leaf_net59),
    .A3(clknet_1_0__leaf_net528),
    .S0(net532),
    .S1(net533),
    .X(net69));
 sky130_fd_sc_hd__mux4_1 c204 (.A0(net840),
    .A1(net1073),
    .A2(clknet_1_0__leaf_net920),
    .A3(net41),
    .S0(net941),
    .S1(net533),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net846),
    .A1(clknet_1_0__leaf_net62),
    .A2(net42),
    .A3(clknet_1_0__leaf_net920),
    .S0(net532),
    .S1(net535),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 c206 (.A0(net46),
    .A1(clknet_1_0__leaf_net62),
    .A2(net532),
    .A3(net533),
    .S0(net535),
    .S1(net536),
    .X(net72));
 sky130_fd_sc_hd__mux4_2 c207 (.A0(net845),
    .A1(net513),
    .A2(net532),
    .A3(net535),
    .S0(net536),
    .S1(net537),
    .X(net925));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(clknet_1_1__leaf_net882),
    .A1(net816),
    .A2(net530),
    .A3(net531),
    .S0(net929),
    .S1(net535),
    .X(net73));
 sky130_fd_sc_hd__mux4_2 c209 (.A0(net849),
    .A1(clknet_1_1__leaf_net73),
    .A2(net925),
    .A3(clknet_1_0__leaf_net62),
    .S0(net535),
    .S1(net537),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 c210 (.A0(net837),
    .A1(net866),
    .A2(net834),
    .A3(net827),
    .S0(net843),
    .S1(clknet_1_0__leaf_net898),
    .X(net904));
 sky130_fd_sc_hd__mux4_1 c211 (.A0(net941),
    .A1(net926),
    .A2(net1067),
    .A3(net865),
    .S0(clknet_1_0__leaf_net57),
    .S1(net48),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(clknet_1_0__leaf_net75),
    .A1(net48),
    .A2(net1019),
    .A3(net1),
    .S0(net943),
    .S1(net929),
    .X(net76));
 sky130_fd_sc_hd__mux4_2 c213 (.A0(net788),
    .A1(net834),
    .A2(net530),
    .A3(net929),
    .S0(net930),
    .S1(net539),
    .X(net876));
 sky130_fd_sc_hd__mux4_2 c214 (.A0(net1),
    .A1(net860),
    .A2(net866),
    .A3(net972),
    .S0(net813),
    .S1(net941),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c215 (.A0(net48),
    .A1(net1068),
    .A2(net859),
    .A3(net784),
    .S0(net800),
    .S1(net910),
    .X(net889));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net994),
    .A1(net876),
    .A2(net839),
    .A3(clknet_1_0__leaf_net57),
    .S0(net949),
    .S1(net813),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_0__leaf_net73),
    .A1(net813),
    .A2(net77),
    .A3(clknet_1_0__leaf_net916),
    .S0(net834),
    .S1(net906),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net1018),
    .A1(net830),
    .A2(net50),
    .A3(clknet_1_0__leaf_net931),
    .S0(net538),
    .S1(net540),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 c219 (.A0(net865),
    .A1(net1067),
    .A2(net944),
    .A3(net850),
    .S0(net791),
    .S1(net1065),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net1006),
    .A1(net986),
    .A2(net943),
    .A3(net810),
    .S0(clknet_1_0__leaf_net904),
    .S1(net541),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 c221 (.A0(net851),
    .A1(net816),
    .A2(clknet_1_0__leaf_net904),
    .A3(net1018),
    .S0(net1006),
    .S1(clknet_1_0__leaf_net528),
    .X(net885));
 sky130_fd_sc_hd__mux4_1 c222 (.A0(clknet_1_1__leaf_net75),
    .A1(net941),
    .A2(clknet_1_0__leaf_net885),
    .A3(net925),
    .S0(net77),
    .S1(net541),
    .X(net83));
 sky130_fd_sc_hd__mux4_2 c223 (.A0(net949),
    .A1(net1075),
    .A2(net0),
    .A3(net1018),
    .S0(net541),
    .S1(net914),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 c224 (.A0(net50),
    .A1(net1049),
    .A2(net1015),
    .A3(net1019),
    .S0(net831),
    .S1(net788),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c225 (.A0(net820),
    .A1(net861),
    .A2(net986),
    .A3(clknet_1_0__leaf_net78),
    .S0(clknet_1_0__leaf_net528),
    .S1(net887),
    .X(net923));
 sky130_fd_sc_hd__mux4_1 c226 (.A0(net784),
    .A1(net850),
    .A2(net1067),
    .A3(net889),
    .S0(net933),
    .S1(net887),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 c227 (.A0(net795),
    .A1(net84),
    .A2(clknet_1_1__leaf_net923),
    .A3(net2),
    .S0(net930),
    .S1(net887),
    .X(net87));
 sky130_fd_sc_hd__mux4_2 c228 (.A0(net84),
    .A1(net809),
    .A2(net86),
    .A3(net951),
    .S0(net1008),
    .S1(net930),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c229 (.A0(net88),
    .A1(clknet_1_0__leaf_net923),
    .A2(net856),
    .A3(clknet_1_0__leaf_net59),
    .S0(net872),
    .S1(net887),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net868),
    .A1(net88),
    .A2(net810),
    .A3(net941),
    .S0(net914),
    .S1(clknet_1_0__leaf_net542),
    .X(net881));
 sky130_fd_sc_hd__a41o_1 c252 (.A1(net1000),
    .A2(net1050),
    .A3(net958),
    .A4(net965),
    .B1(net996),
    .X(net875));
 sky130_fd_sc_hd__a41o_2 c253 (.A1(net955),
    .A2(net1054),
    .A3(net959),
    .A4(net1011),
    .B1(net1071),
    .X(net90));
 sky130_fd_sc_hd__a41o_2 c254 (.A1(net1011),
    .A2(net814),
    .A3(net954),
    .A4(net1056),
    .B1(net1019),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(net1056),
    .A1(net1018),
    .A2(net954),
    .A3(net1002),
    .S0(net983),
    .S1(net962),
    .X(net92));
 sky130_fd_sc_hd__a41o_2 c256 (.A1(net979),
    .A2(net21),
    .A3(net994),
    .A4(net955),
    .B1(net952),
    .X(net93));
 sky130_fd_sc_hd__a41o_2 c257 (.A1(net1015),
    .A2(net1055),
    .A3(net954),
    .A4(net952),
    .B1(net93),
    .X(net94));
 sky130_fd_sc_hd__sdfbbn_2 c258 (.CLK_N(clknet_leaf_8_clk),
    .D(net20),
    .RESET_B(net90),
    .SCD(net94),
    .SCE(net1055),
    .SET_B(net955),
    .Q(net900),
    .Q_N(net95));
 sky130_fd_sc_hd__a41o_4 c259 (.A1(net900),
    .A2(net1024),
    .A3(net955),
    .A4(net1055),
    .B1(net1056),
    .X(net96));
 sky130_fd_sc_hd__mux4_2 c260 (.A0(net96),
    .A1(net90),
    .A2(net93),
    .A3(net955),
    .S0(net1057),
    .S1(net952),
    .X(net97));
 sky130_fd_sc_hd__a41o_2 c261 (.A1(net1019),
    .A2(net1011),
    .A3(net91),
    .A4(net954),
    .B1(net1055),
    .X(net98));
 sky130_fd_sc_hd__sdfbbn_1 c262 (.CLK_N(clknet_leaf_9_clk),
    .D(net93),
    .RESET_B(net94),
    .SCD(net96),
    .SCE(net97),
    .SET_B(net954),
    .Q(net100),
    .Q_N(net99));
 sky130_fd_sc_hd__sdfbbp_1 c263 (.CLK(clknet_leaf_9_clk),
    .D(net1054),
    .RESET_B(net94),
    .SCD(net98),
    .SCE(net1074),
    .SET_B(net954),
    .Q(net102),
    .Q_N(net101));
 sky130_fd_sc_hd__mux4_2 c264 (.A0(net100),
    .A1(net93),
    .A2(net1018),
    .A3(net954),
    .S0(net1057),
    .S1(net101),
    .X(net103));
 sky130_fd_sc_hd__mux4_1 c265 (.A0(net97),
    .A1(net100),
    .A2(net814),
    .A3(net954),
    .S0(net1056),
    .S1(net1071),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 c266 (.A0(net997),
    .A1(net102),
    .A2(net99),
    .A3(net1058),
    .S0(net954),
    .S1(net97),
    .X(net105));
 sky130_fd_sc_hd__mux4_1 c267 (.A0(net94),
    .A1(net900),
    .A2(net1014),
    .A3(net99),
    .S0(net955),
    .S1(net101),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c268 (.A0(net90),
    .A1(net97),
    .A2(net103),
    .A3(net94),
    .S0(net962),
    .S1(net545),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c269 (.A0(net1072),
    .A1(net93),
    .A2(net103),
    .A3(net96),
    .S0(net95),
    .S1(net546),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 c270 (.A0(net98),
    .A1(net103),
    .A2(net1075),
    .A3(net101),
    .S0(clknet_1_0__leaf_net543),
    .S1(net547),
    .X(net109));
 sky130_fd_sc_hd__mux4_2 c271 (.A0(net91),
    .A1(net98),
    .A2(net101),
    .A3(net1101),
    .S0(net547),
    .S1(net548),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(net110),
    .A1(net93),
    .A2(net96),
    .A3(clknet_1_1__leaf_net543),
    .S0(net547),
    .S1(net549),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 c273 (.A0(net1024),
    .A1(net1069),
    .A2(net1000),
    .A3(net1006),
    .S0(net952),
    .S1(clknet_1_1__leaf_net544),
    .X(net112));
 sky130_fd_sc_hd__mux4_2 c274 (.A0(net783),
    .A1(net800),
    .A2(net791),
    .A3(net1019),
    .S0(net946),
    .S1(net525),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 c275 (.A0(clknet_1_1__leaf_net112),
    .A1(net27),
    .A2(net962),
    .A3(net965),
    .S0(net952),
    .S1(net1071),
    .X(net114));
 sky130_fd_sc_hd__a41o_1 c276 (.A1(net926),
    .A2(clknet_1_0__leaf_net114),
    .A3(net1010),
    .A4(net9),
    .B1(net525),
    .X(net115));
 sky130_fd_sc_hd__a41o_1 c277 (.A1(clknet_1_0__leaf_net114),
    .A2(net98),
    .A3(net789),
    .A4(net512),
    .B1(net523),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 c278 (.A0(net1073),
    .A1(net99),
    .A2(net33),
    .A3(net95),
    .S0(net990),
    .S1(net980),
    .X(net117));
 sky130_fd_sc_hd__mux4_1 c279 (.A0(net793),
    .A1(net4),
    .A2(net799),
    .A3(net972),
    .S0(clknet_1_1__leaf_net116),
    .S1(clknet_1_1__leaf_net544),
    .X(net883));
 sky130_fd_sc_hd__mux4_1 c280 (.A0(net789),
    .A1(net1072),
    .A2(clknet_1_1__leaf_net883),
    .A3(net525),
    .S0(net547),
    .S1(net551),
    .X(net118));
 sky130_fd_sc_hd__mux4_1 c281 (.A0(net999),
    .A1(net113),
    .A2(net979),
    .A3(net19),
    .S0(net798),
    .S1(clknet_1_1__leaf_net883),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net798),
    .A1(net949),
    .A2(clknet_1_1__leaf_net883),
    .A3(net548),
    .S0(net551),
    .S1(net552),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 c283 (.A0(clknet_1_1__leaf_net883),
    .A1(net952),
    .A2(net990),
    .A3(clknet_1_1__leaf_net112),
    .S0(net999),
    .S1(net553),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 c284 (.A0(net793),
    .A1(clknet_1_0__leaf_net116),
    .A2(net779),
    .A3(net997),
    .S0(net512),
    .S1(net553),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net1035),
    .A1(clknet_1_1__leaf_net115),
    .A2(clknet_1_1__leaf_net116),
    .A3(net103),
    .S0(net949),
    .S1(net519),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 c286 (.A0(net800),
    .A1(clknet_1_1__leaf_net114),
    .A2(clknet_1_1__leaf_net883),
    .A3(net1073),
    .S0(net551),
    .S1(net553),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 c287 (.A0(net990),
    .A1(clknet_1_1__leaf_net883),
    .A2(net526),
    .A3(clknet_1_0__leaf_net543),
    .S0(net554),
    .S1(net555),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(clknet_1_1__leaf_net116),
    .A1(net943),
    .A2(net991),
    .A3(clknet_1_1__leaf_net883),
    .S0(net552),
    .S1(net557),
    .X(net126));
 sky130_fd_sc_hd__mux4_2 c289 (.A0(net93),
    .A1(net1022),
    .A2(net1086),
    .A3(net553),
    .S0(net559),
    .S1(net560),
    .X(net919));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net103),
    .A1(net783),
    .A2(net919),
    .A3(net790),
    .S0(net555),
    .S1(net559),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 c291 (.A0(net798),
    .A1(clknet_1_0__leaf_net111),
    .A2(net547),
    .A3(net556),
    .S0(net557),
    .S1(net561),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 c292 (.A0(clknet_1_1__leaf_net115),
    .A1(clknet_1_1__leaf_net883),
    .A2(net919),
    .A3(net553),
    .S0(net560),
    .S1(clknet_1_0__leaf_net562),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 c293 (.A0(net33),
    .A1(net793),
    .A2(clknet_1_1__leaf_net883),
    .A3(net519),
    .S0(net559),
    .S1(net561),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 c294 (.A0(clknet_1_0__leaf_net54),
    .A1(clknet_1_1__leaf_net57),
    .A2(net821),
    .A3(net804),
    .S0(net816),
    .S1(clknet_1_0__leaf_net544),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c295 (.A0(net828),
    .A1(clknet_1_0__leaf_net131),
    .A2(net823),
    .A3(net20),
    .S0(clknet_1_0__leaf_net529),
    .S1(net559),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c296 (.A0(net822),
    .A1(clknet_1_0__leaf_net114),
    .A2(net950),
    .A3(net999),
    .S0(net1015),
    .S1(clknet_1_1__leaf_net529),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 c297 (.A0(clknet_1_0__leaf_net116),
    .A1(clknet_1_1__leaf_net133),
    .A2(net919),
    .A3(net18),
    .S0(net1012),
    .S1(net980),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 c298 (.A0(net23),
    .A1(clknet_1_1__leaf_net882),
    .A2(net1069),
    .A3(net957),
    .S0(clknet_1_0__leaf_net132),
    .S1(net526),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(clknet_1_1__leaf_net133),
    .A1(net1054),
    .A2(net1071),
    .A3(net826),
    .S0(net31),
    .S1(clknet_1_0__leaf_net562),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 c300 (.A0(net821),
    .A1(clknet_1_1__leaf_net54),
    .A2(net1014),
    .A3(net814),
    .S0(net961),
    .S1(net798),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 c301 (.A0(clknet_1_0__leaf_net116),
    .A1(clknet_1_1__leaf_net883),
    .A2(net52),
    .A3(net551),
    .S0(clknet_1_0__leaf_net563),
    .S1(net564),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 c302 (.A0(clknet_1_0__leaf_net132),
    .A1(net984),
    .A2(net822),
    .A3(net46),
    .S0(net41),
    .S1(net526),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 c303 (.A0(net828),
    .A1(net979),
    .A2(clknet_1_1__leaf_net136),
    .A3(net1012),
    .S1(net566),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net793),
    .A1(clknet_1_1__leaf_net137),
    .A2(clknet_1_1__leaf_net133),
    .A3(net948),
    .S0(net982),
    .S1(net567),
    .X(net899));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net508),
    .A1(net511),
    .A2(net552),
    .A3(clknet_1_1__leaf_net563),
    .S0(net564),
    .S1(net567),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net46),
    .A1(net1003),
    .A2(net980),
    .A3(net559),
    .S0(clknet_1_0__leaf_net563),
    .S1(net566),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(clknet_1_0__leaf_net137),
    .A1(net98),
    .A2(clknet_1_1__leaf_net132),
    .A3(clknet_1_0__leaf_net141),
    .S0(net564),
    .S1(net566),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net1023),
    .A1(clknet_1_1__leaf_net132),
    .A2(clknet_1_0__leaf_net137),
    .A3(net511),
    .S0(clknet_1_0__leaf_net563),
    .S1(net568),
    .X(net144));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net1023),
    .A1(clknet_1_1__leaf_net899),
    .A2(clknet_1_1__leaf_net136),
    .A3(clknet_1_0__leaf_net142),
    .S0(net553),
    .S1(net568),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(clknet_1_0__leaf_net136),
    .A1(clknet_1_0__leaf_net133),
    .A2(clknet_1_1__leaf_net899),
    .A3(net511),
    .S0(clknet_1_0__leaf_net563),
    .S1(net570),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 c311 (.A0(clknet_1_0__leaf_net141),
    .A1(clknet_1_0__leaf_net529),
    .A2(clknet_1_1__leaf_net908),
    .A3(net566),
    .S0(net570),
    .S1(net571),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(clknet_1_0__leaf_net147),
    .A1(net821),
    .A2(net1067),
    .A3(clknet_1_0__leaf_net563),
    .S0(net565),
    .S1(net571),
    .X(net884));
 sky130_fd_sc_hd__mux4_1 c313 (.A0(net31),
    .A1(clknet_1_1__leaf_net147),
    .A2(net1030),
    .A3(clknet_1_0__leaf_net563),
    .S0(net570),
    .S1(net571),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 c314 (.A0(net1075),
    .A1(clknet_1_1__leaf_net112),
    .A2(clknet_1_0__leaf_net148),
    .A3(net907),
    .S0(net570),
    .S1(net571),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 c315 (.A0(net823),
    .A1(net1034),
    .A2(net95),
    .A3(net973),
    .S0(net94),
    .S1(clknet_1_1__leaf_net64),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(clknet_1_0__leaf_net142),
    .A1(net1018),
    .A2(net814),
    .A3(net961),
    .S0(net507),
    .S1(net535),
    .X(net893));
 sky130_fd_sc_hd__mux4_1 c317 (.A0(clknet_1_1__leaf_net899),
    .A1(net52),
    .A2(net828),
    .A3(net838),
    .S0(net1071),
    .S1(net507),
    .X(net151));
 sky130_fd_sc_hd__mux4_2 c318 (.A0(net1054),
    .A1(net809),
    .A2(net967),
    .A3(net521),
    .S0(net531),
    .S1(net552),
    .X(net913));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net94),
    .A1(clknet_1_0__leaf_net883),
    .A2(net919),
    .A3(net835),
    .S0(net913),
    .S1(net535),
    .X(net152));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net1018),
    .A1(net835),
    .A2(net838),
    .A3(net1002),
    .S0(clknet_1_1__leaf_net528),
    .S1(net569),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(clknet_1_1__leaf_net153),
    .A1(clknet_1_0__leaf_net133),
    .A2(clknet_1_0__leaf_net122),
    .A3(net997),
    .S0(net972),
    .S1(net982),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(net41),
    .A1(net972),
    .A2(net817),
    .A3(clknet_1_1__leaf_net893),
    .S0(net577),
    .S1(net578),
    .X(net155));
 sky130_fd_sc_hd__mux4_2 c323 (.A0(clknet_1_0__leaf_net147),
    .A1(net46),
    .A2(net807),
    .A3(clknet_1_1__leaf_net59),
    .S0(net571),
    .S1(net576),
    .X(net156));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(net835),
    .A1(clknet_1_1__leaf_net920),
    .A2(net999),
    .A3(net813),
    .S0(net1060),
    .S1(net578),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 c325 (.A0(net828),
    .A1(net841),
    .A2(net809),
    .A3(net948),
    .S0(clknet_1_1__leaf_net528),
    .S1(net576),
    .X(net158));
 sky130_fd_sc_hd__mux4_2 c326 (.A0(clknet_1_0__leaf_net156),
    .A1(net1074),
    .A2(net1003),
    .A3(net951),
    .S0(net578),
    .S1(net911),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(clknet_1_0__leaf_net153),
    .A1(net941),
    .A2(net1011),
    .A3(net913),
    .S0(net573),
    .S1(net574),
    .X(net160));
 sky130_fd_sc_hd__sdfbbn_1 c328 (.CLK_N(clknet_leaf_42_clk),
    .D(net826),
    .RESET_B(net1104),
    .SCD(net943),
    .SCE(net517),
    .SET_B(net1064),
    .Q(net162),
    .Q_N(net161));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net136),
    .A1(clknet_1_0__leaf_net64),
    .A2(clknet_1_0__leaf_net159),
    .A3(net906),
    .S0(net535),
    .S1(net578),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net787),
    .A1(net816),
    .A2(net804),
    .A3(net1081),
    .S0(net1006),
    .S1(net577),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c331 (.A0(clknet_1_1__leaf_net156),
    .A1(net972),
    .A2(net1002),
    .A3(net941),
    .S0(net537),
    .S1(clknet_1_0__leaf_net580),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net838),
    .A1(clknet_1_0__leaf_net165),
    .A2(net906),
    .A3(clknet_1_0__leaf_net883),
    .S0(net574),
    .S1(net578),
    .X(net166));
 sky130_fd_sc_hd__mux4_2 c333 (.A0(clknet_1_1__leaf_net153),
    .A1(clknet_1_0__leaf_net159),
    .A2(net835),
    .S0(net521),
    .S1(net578),
    .X(net918));
 sky130_fd_sc_hd__mux4_1 c334 (.A0(clknet_1_0__leaf_net64),
    .A1(clknet_1_0__leaf_net165),
    .A2(net833),
    .A3(net161),
    .S0(clknet_1_1__leaf_net893),
    .S1(clknet_1_0__leaf_net580),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 c335 (.A0(clknet_1_0__leaf_net165),
    .A1(net1054),
    .A2(clknet_1_1__leaf_net159),
    .A3(clknet_1_1__leaf_net918),
    .S0(clknet_1_1__leaf_net580),
    .S1(clknet_1_1__leaf_net902),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(net97),
    .A1(net856),
    .A2(net88),
    .A3(net853),
    .S0(net984),
    .S1(net854),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 c337 (.A0(net797),
    .A1(net854),
    .A2(net814),
    .A3(net1018),
    .S0(clknet_1_0__leaf_net883),
    .S1(clknet_1_0__leaf_net115),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 c338 (.A0(clknet_1_0__leaf_net83),
    .A1(net853),
    .A2(clknet_1_0__leaf_net62),
    .A3(net854),
    .S0(net561),
    .S1(net909),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net0),
    .A1(net844),
    .A2(net862),
    .A3(net103),
    .S0(net910),
    .S1(net584),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_0__leaf_net160),
    .A1(net0),
    .A2(net852),
    .A3(net97),
    .S0(net913),
    .S1(clknet_1_0__leaf_net528),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(clknet_1_0__leaf_net122),
    .A1(clknet_1_0__leaf_net153),
    .A2(net913),
    .A3(net941),
    .S0(net1075),
    .S1(net584),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c342 (.A0(net859),
    .A1(net1051),
    .A2(net926),
    .A3(clknet_1_0__leaf_net882),
    .S0(net565),
    .S1(net586),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net790),
    .A1(clknet_1_1__leaf_net160),
    .A2(net86),
    .A3(net1010),
    .S0(net579),
    .S1(net584),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(net88),
    .A1(net961),
    .A2(net841),
    .A3(net864),
    .S0(clknet_1_1__leaf_net908),
    .S1(net587),
    .X(net178));
 sky130_fd_sc_hd__mux4_2 c345 (.A0(clknet_1_0__leaf_net61),
    .A1(net876),
    .A2(net841),
    .A3(net800),
    .S0(clknet_1_0__leaf_net178),
    .S1(net855),
    .X(net870));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net86),
    .A1(net926),
    .A2(net854),
    .A3(clknet_1_1__leaf_net904),
    .S0(net534),
    .S1(net586),
    .X(net901));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net949),
    .A1(clknet_1_0__leaf_net899),
    .A2(net859),
    .A3(net855),
    .S0(net585),
    .S1(net586),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(clknet_1_1__leaf_net899),
    .A1(net941),
    .A2(clknet_1_0__leaf_net178),
    .A3(net161),
    .S0(net570),
    .S1(net586),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net77),
    .A1(net1003),
    .A2(net534),
    .A3(net582),
    .S0(net909),
    .S1(net589),
    .X(net917));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(net841),
    .A1(clknet_1_0__leaf_net870),
    .A2(net88),
    .A3(net579),
    .S0(clknet_1_0__leaf_net902),
    .S1(net586),
    .X(net181));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net103),
    .A1(clknet_1_1__leaf_net83),
    .A2(net889),
    .A3(net515),
    .S0(net911),
    .S1(net590),
    .X(net182));
 sky130_fd_sc_hd__mux4_1 c352 (.A0(clknet_1_0__leaf_net57),
    .A1(clknet_1_0__leaf_net870),
    .A2(clknet_1_0__leaf_net908),
    .A3(net573),
    .S0(net590),
    .S1(net593),
    .X(net183));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(net1067),
    .A1(clknet_1_0__leaf_net178),
    .A2(net162),
    .A3(net909),
    .S0(net586),
    .S1(net591),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 c354 (.A0(clknet_1_1__leaf_net920),
    .A1(clknet_1_0__leaf_net884),
    .A2(net97),
    .A3(net516),
    .S0(net589),
    .S1(net592),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net176),
    .A1(net1041),
    .A2(clknet_1_0__leaf_net918),
    .A3(net571),
    .S0(net591),
    .S1(net594),
    .X(net903));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(clknet_1_0__leaf_net870),
    .A1(net866),
    .A2(clknet_1_0__leaf_net178),
    .A3(net905),
    .S0(net591),
    .S1(net594),
    .X(net186));
 sky130_fd_sc_hd__sdfbbn_2 c378 (.CLK_N(clknet_leaf_12_clk),
    .D(net102),
    .RESET_B(net167),
    .SCD(clknet_1_1__leaf_net111),
    .SCE(net1059),
    .SET_B(net1032),
    .Q(net188),
    .Q_N(net187));
 sky130_fd_sc_hd__a41o_2 c379 (.A1(net984),
    .A2(net964),
    .A3(net952),
    .A4(net951),
    .B1(net167),
    .X(net189));
 sky130_fd_sc_hd__a41o_4 c380 (.A1(net188),
    .A2(net167),
    .A3(net772),
    .A4(net1000),
    .B1(net189),
    .X(net871));
 sky130_fd_sc_hd__a41o_2 c381 (.A1(net167),
    .A2(net871),
    .A3(net95),
    .A4(net992),
    .B1(net954),
    .X(net190));
 sky130_fd_sc_hd__a41o_1 c382 (.A1(net964),
    .A2(net1072),
    .A3(net190),
    .A4(net91),
    .B1(net101),
    .X(net191));
 sky130_fd_sc_hd__a41o_1 c383 (.A1(net953),
    .A2(net871),
    .A3(net96),
    .A4(net992),
    .B1(net549),
    .X(net192));
 sky130_fd_sc_hd__mux4_2 c384 (.A0(net1059),
    .A1(net1072),
    .A2(net11),
    .A3(net991),
    .S0(net545),
    .S1(net980),
    .X(net873));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(net989),
    .A1(clknet_1_1__leaf_net111),
    .A2(net190),
    .A3(net192),
    .S0(net992),
    .S1(clknet_1_1__leaf_net543),
    .X(net193));
 sky130_fd_sc_hd__a41o_1 c386 (.A1(net873),
    .A2(net192),
    .A3(net190),
    .A4(net871),
    .B1(clknet_1_1__leaf_net543),
    .X(net897));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net994),
    .A1(net102),
    .A2(net167),
    .A3(clknet_1_1__leaf_net897),
    .S0(net192),
    .S1(net503),
    .X(net194));
 sky130_fd_sc_hd__sdfbbp_1 c388 (.CLK(clknet_leaf_10_clk),
    .D(net1072),
    .RESET_B(clknet_1_1__leaf_net111),
    .SCD(net945),
    .SCE(clknet_1_0__leaf_net897),
    .SET_B(clknet_1_1__leaf_net544),
    .Q(net196),
    .Q_N(net195));
 sky130_fd_sc_hd__a41o_1 c389 (.A1(net190),
    .A2(net196),
    .A3(net945),
    .A4(net91),
    .B1(net503),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net942),
    .A1(clknet_1_1__leaf_net194),
    .A2(net195),
    .A3(net955),
    .S0(net989),
    .S1(net546),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(net196),
    .A1(net942),
    .A2(clknet_1_1__leaf_net897),
    .A3(net503),
    .S0(net545),
    .S1(clknet_1_0__leaf_net596),
    .X(net199));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net167),
    .A1(clknet_1_0__leaf_net897),
    .A2(net942),
    .A3(net952),
    .S0(net195),
    .S1(net980),
    .X(net200));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net196),
    .A1(net1015),
    .A2(net942),
    .A3(clknet_1_0__leaf_net596),
    .S0(clknet_1_1__leaf_net597),
    .S1(clknet_1_0__leaf_net598),
    .X(net201));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(clknet_1_1__leaf_net194),
    .A1(net921),
    .A2(net195),
    .A3(net549),
    .S0(clknet_1_1__leaf_net597),
    .S1(clknet_1_0__leaf_net598),
    .X(net202));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(net871),
    .A1(net192),
    .A2(clknet_1_0__leaf_net194),
    .A3(clknet_1_0__leaf_net598),
    .S0(net600),
    .S1(net601),
    .X(net203));
 sky130_fd_sc_hd__mux4_1 c396 (.A0(net956),
    .A1(net190),
    .A2(net960),
    .A3(clknet_1_0__leaf_net596),
    .S0(net600),
    .S1(net604),
    .X(net204));
 sky130_fd_sc_hd__mux4_1 c397 (.A0(clknet_1_1__leaf_net897),
    .A1(net942),
    .A2(clknet_1_1__leaf_net204),
    .A3(net100),
    .S0(clknet_1_1__leaf_net598),
    .S1(net599),
    .X(net205));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net942),
    .A1(net980),
    .A2(clknet_1_1__leaf_net597),
    .A3(net602),
    .S0(net603),
    .S1(net605),
    .X(net206));
 sky130_fd_sc_hd__mux4_1 c399 (.A0(net1006),
    .A1(net1046),
    .A2(net519),
    .A3(net524),
    .S0(clknet_1_0__leaf_net543),
    .S1(net555),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 c400 (.A0(net1000),
    .A1(net797),
    .A2(net99),
    .A3(net12),
    .S0(net1002),
    .S1(net560),
    .X(net208));
 sky130_fd_sc_hd__mux4_1 c401 (.A0(net100),
    .A1(net33),
    .A2(clknet_1_0__leaf_net207),
    .A3(clknet_1_0__leaf_net194),
    .S0(net1006),
    .S1(clknet_1_1__leaf_net883),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 c402 (.A0(net797),
    .A1(net943),
    .A2(net946),
    .A3(net942),
    .S0(clknet_1_1__leaf_net883),
    .S1(net519),
    .X(net210));
 sky130_fd_sc_hd__mux4_2 c403 (.A0(net796),
    .A1(net208),
    .A2(net98),
    .A3(net1031),
    .S0(net959),
    .S1(net606),
    .X(net211));
 sky130_fd_sc_hd__mux4_1 c404 (.A0(net783),
    .A1(net211),
    .A2(net942),
    .A3(net802),
    .S0(net551),
    .S1(net606),
    .X(net212));
 sky130_fd_sc_hd__mux4_1 c405 (.A0(net211),
    .A1(net991),
    .A2(clknet_1_0__leaf_net111),
    .A3(net919),
    .S0(net1001),
    .S1(clknet_1_0__leaf_net596),
    .X(net213));
 sky130_fd_sc_hd__mux4_1 c406 (.A0(net1006),
    .A1(clknet_1_0__leaf_net111),
    .A2(net1001),
    .A3(net554),
    .S0(clknet_1_0__leaf_net562),
    .S1(net608),
    .X(net214));
 sky130_fd_sc_hd__mux4_2 c407 (.A0(net952),
    .A1(net915),
    .A2(net525),
    .A3(net560),
    .S0(net608),
    .S1(net878),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c408 (.A0(net113),
    .A1(net215),
    .A2(net197),
    .A3(net991),
    .S0(net512),
    .S1(net606),
    .X(net216));
 sky130_fd_sc_hd__mux4_1 c409 (.A0(clknet_1_0__leaf_net111),
    .A1(net90),
    .A2(net797),
    .A3(net96),
    .S0(net606),
    .S1(net608),
    .X(net217));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net21),
    .A1(net208),
    .A2(net796),
    .A3(net886),
    .S0(net606),
    .S1(net613),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c411 (.A0(clknet_1_0__leaf_net194),
    .A1(net873),
    .A2(net991),
    .A3(net785),
    .S0(net218),
    .S1(net548),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c412 (.A0(net1022),
    .A1(clknet_1_0__leaf_net207),
    .A2(net785),
    .A3(net218),
    .S0(net802),
    .S1(net980),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c413 (.A0(clknet_1_1__leaf_net220),
    .A1(net952),
    .A2(net980),
    .A3(net606),
    .S0(net608),
    .S1(net614),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net945),
    .A1(net101),
    .A2(clknet_1_1__leaf_net543),
    .A3(net549),
    .S0(net611),
    .S1(net615),
    .X(net222));
 sky130_fd_sc_hd__mux4_1 c415 (.A0(net1038),
    .A1(clknet_1_1__leaf_net220),
    .A2(net524),
    .A3(net607),
    .S0(net609),
    .S1(net613),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(clknet_1_0__leaf_net207),
    .A1(clknet_1_0__leaf_net222),
    .A2(net988),
    .A3(clknet_1_1__leaf_net220),
    .S0(net614),
    .S1(clknet_1_0__leaf_net616),
    .X(net224));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net1014),
    .A1(net189),
    .A2(clknet_1_1__leaf_net220),
    .A3(net556),
    .S0(net615),
    .S1(clknet_1_0__leaf_net616),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c418 (.A0(net873),
    .A1(net218),
    .A2(net615),
    .A3(clknet_1_1__leaf_net616),
    .S0(clknet_1_0__leaf_net617),
    .S1(clknet_1_1__leaf_net618),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net21),
    .A1(clknet_1_0__leaf_net222),
    .A2(clknet_1_0__leaf_net226),
    .A3(clknet_1_1__leaf_net220),
    .S0(net614),
    .S1(clknet_1_0__leaf_net617),
    .X(net227));
 sky130_fd_sc_hd__mux4_1 c420 (.A0(net98),
    .A1(clknet_1_1__leaf_net122),
    .A2(net40),
    .A3(clknet_1_1__leaf_net884),
    .S0(net1037),
    .S1(net606),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c421 (.A0(clknet_1_0__leaf_net142),
    .A1(net826),
    .A2(net511),
    .A3(net527),
    .S0(net569),
    .S1(net614),
    .X(net229));
 sky130_fd_sc_hd__mux4_2 c422 (.A0(net1034),
    .A1(net1009),
    .A2(net783),
    .A3(net43),
    .S0(net522),
    .S1(net605),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 c423 (.A0(clknet_1_0__leaf_net131),
    .A1(clknet_1_0__leaf_net148),
    .A2(clknet_1_0__leaf_net229),
    .A3(net90),
    .S0(net1034),
    .S1(net611),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c424 (.A0(net797),
    .A1(net215),
    .A2(net919),
    .A3(net1003),
    .S0(net1008),
    .S1(net1032),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c425 (.A0(net783),
    .A1(net991),
    .A2(clknet_1_0__leaf_net229),
    .A3(net567),
    .S0(net569),
    .S1(net622),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c426 (.A0(net1037),
    .A1(clknet_1_1__leaf_net141),
    .A2(net1003),
    .A3(net999),
    .S0(net211),
    .S1(net621),
    .X(net234));
 sky130_fd_sc_hd__mux4_2 c427 (.A0(net90),
    .A1(net945),
    .A2(net946),
    .A3(net607),
    .S0(net613),
    .S1(net621),
    .X(net928));
 sky130_fd_sc_hd__mux4_1 c428 (.A0(clknet_1_1__leaf_net148),
    .A1(clknet_1_1__leaf_net122),
    .A2(net817),
    .A3(clknet_1_0__leaf_net220),
    .S0(net1029),
    .S1(clknet_1_0__leaf_net597),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c429 (.A0(clknet_1_1__leaf_net141),
    .A1(clknet_1_0__leaf_net226),
    .A2(net797),
    .A3(net1053),
    .S0(clknet_1_1__leaf_net148),
    .S1(net600),
    .X(net236));
 sky130_fd_sc_hd__mux4_1 c430 (.A0(net211),
    .A1(net962),
    .A2(net967),
    .A3(clknet_1_1__leaf_net148),
    .S0(net612),
    .S1(net623),
    .X(net237));
 sky130_fd_sc_hd__mux4_1 c431 (.A0(net945),
    .A1(clknet_1_0__leaf_net883),
    .A2(net919),
    .A3(clknet_1_0__leaf_net897),
    .S0(net511),
    .S1(net626),
    .X(net238));
 sky130_fd_sc_hd__mux4_2 c432 (.A0(net817),
    .A1(net988),
    .A2(net52),
    .A3(net551),
    .S0(net610),
    .S1(net612),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 c433 (.A0(net230),
    .A1(clknet_1_1__leaf_net133),
    .A2(net886),
    .A3(clknet_1_1__leaf_net563),
    .S0(net567),
    .S1(clknet_1_0__leaf_net597),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 c434 (.A0(net1009),
    .A1(net1011),
    .A2(net40),
    .A3(net511),
    .S0(net567),
    .S1(clknet_1_0__leaf_net597),
    .X(net241));
 sky130_fd_sc_hd__mux4_1 c435 (.A0(clknet_1_0__leaf_net241),
    .A1(net37),
    .A2(clknet_1_1__leaf_net229),
    .A3(net819),
    .S0(net613),
    .S1(net622),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net211),
    .A1(clknet_1_0__leaf_net882),
    .A2(net569),
    .A3(net606),
    .S0(net607),
    .S1(net628),
    .X(net243));
 sky130_fd_sc_hd__mux4_1 c437 (.A0(clknet_1_1__leaf_net243),
    .A1(net783),
    .A2(net509),
    .A3(net605),
    .S0(net625),
    .S1(net628),
    .X(net244));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(clknet_1_0__leaf_net241),
    .A1(net90),
    .A2(clknet_1_1__leaf_net240),
    .A3(clknet_1_1__leaf_net243),
    .S0(net606),
    .S1(net629),
    .X(net245));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(clknet_1_0__leaf_net240),
    .A1(clknet_1_1__leaf_net131),
    .A2(net928),
    .A3(net1035),
    .S0(net527),
    .S1(net629),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(clknet_1_1__leaf_net233),
    .A1(net807),
    .A2(clknet_1_1__leaf_net563),
    .A3(net629),
    .S0(net630),
    .S1(net632),
    .X(net247));
 sky130_fd_sc_hd__mux4_1 c441 (.A0(net21),
    .A1(net796),
    .A2(clknet_1_1__leaf_net59),
    .A3(net972),
    .S0(net578),
    .S1(net629),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c442 (.A0(net1032),
    .A1(net1010),
    .A2(clknet_1_0__leaf_net226),
    .A3(net999),
    .S0(net844),
    .S1(net187),
    .X(net249));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net1081),
    .A1(clknet_1_0__leaf_net62),
    .A2(net997),
    .A3(net833),
    .S0(net943),
    .S1(net844),
    .X(net250));
 sky130_fd_sc_hd__mux4_1 c444 (.A0(clknet_1_1__leaf_net159),
    .A1(net188),
    .A2(clknet_1_1__leaf_net243),
    .A3(net1028),
    .S0(net96),
    .S1(net790),
    .X(net251));
 sky130_fd_sc_hd__mux4_1 c445 (.A0(net215),
    .A1(net1034),
    .A2(clknet_1_1__leaf_net122),
    .A3(net967),
    .S0(net808),
    .S1(net1002),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c446 (.A0(clknet_1_1__leaf_net59),
    .A1(clknet_1_1__leaf_net47),
    .A2(net986),
    .A3(net575),
    .S0(net623),
    .S1(net627),
    .X(net253));
 sky130_fd_sc_hd__mux4_1 c447 (.A0(net946),
    .A1(clknet_1_1__leaf_net59),
    .A2(net564),
    .A3(net578),
    .S0(net634),
    .S1(net635),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(clknet_1_0__leaf_net248),
    .A1(net162),
    .A2(clknet_1_0__leaf_net133),
    .A3(net1073),
    .S0(net984),
    .S1(net537),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 c449 (.A0(net1034),
    .A1(net919),
    .A2(clknet_1_1__leaf_net248),
    .A3(net537),
    .S0(net569),
    .S1(net575),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net839),
    .A1(net1077),
    .A2(clknet_1_0__leaf_net233),
    .A3(net21),
    .S0(net634),
    .S1(clknet_1_1__leaf_net637),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 c451 (.A0(clknet_1_1__leaf_net898),
    .A1(net578),
    .A2(clknet_1_1__leaf_net618),
    .A3(net627),
    .S0(net636),
    .S1(clknet_1_1__leaf_net637),
    .X(net258));
 sky130_fd_sc_hd__mux4_1 c452 (.A0(clknet_1_0__leaf_net255),
    .A1(clknet_1_0__leaf_net257),
    .A2(net164),
    .A3(net841),
    .S0(net839),
    .S1(clknet_1_0__leaf_net637),
    .X(net259));
 sky130_fd_sc_hd__mux4_1 c453 (.A0(clknet_1_0__leaf_net258),
    .A1(net972),
    .A2(net841),
    .A3(net994),
    .S0(net630),
    .S1(clknet_1_1__leaf_net637),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 c454 (.A0(net817),
    .A1(net1019),
    .A2(clknet_1_1__leaf_net258),
    .A3(clknet_1_1__leaf_net253),
    .S0(clknet_1_1__leaf_net260),
    .S1(net520),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 c455 (.A0(clknet_1_0__leaf_net260),
    .A1(net997),
    .A2(clknet_1_1__leaf_net255),
    .A3(net1008),
    .S0(net578),
    .S1(clknet_1_0__leaf_net581),
    .X(net262));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(clknet_1_1__leaf_net254),
    .A1(clknet_1_1__leaf_net261),
    .A2(net531),
    .A3(net558),
    .S0(clknet_1_0__leaf_net581),
    .S1(clknet_1_1__leaf_net638),
    .X(net263));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net833),
    .A1(clknet_1_0__leaf_net122),
    .A2(net230),
    .A3(net558),
    .S0(clknet_1_0__leaf_net637),
    .S1(net639),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net164),
    .A1(clknet_1_0__leaf_net257),
    .A2(net635),
    .A3(clknet_1_0__leaf_net637),
    .S0(net639),
    .S1(net641),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(clknet_1_0__leaf_net261),
    .A1(clknet_1_0__leaf_net254),
    .A2(net21),
    .A3(clknet_1_1__leaf_net62),
    .S0(clknet_1_1__leaf_net637),
    .S1(net640),
    .X(net266));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(clknet_1_0__leaf_net257),
    .A1(net1010),
    .A2(clknet_1_1__leaf_net898),
    .A3(clknet_1_0__leaf_net637),
    .S0(clknet_1_0__leaf_net638),
    .S1(net639),
    .X(net267));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(clknet_1_1__leaf_net257),
    .A1(net520),
    .A2(net575),
    .A3(clknet_1_0__leaf_net638),
    .S0(net642),
    .S1(net645),
    .X(net268));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net1041),
    .A1(net943),
    .A2(clknet_1_0__leaf_net112),
    .A3(clknet_1_1__leaf_net47),
    .S0(clknet_1_1__leaf_net885),
    .S1(net864),
    .X(net269));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net1053),
    .A1(net852),
    .A2(net864),
    .A3(net973),
    .S0(clknet_1_1__leaf_net542),
    .S1(net589),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net854),
    .A1(net1041),
    .A2(net864),
    .A3(clknet_1_1__leaf_net870),
    .S0(clknet_1_0__leaf_net899),
    .S1(net586),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net96),
    .A1(net816),
    .A2(clknet_1_0__leaf_net897),
    .A3(net1010),
    .S0(net514),
    .S1(net589),
    .X(net272));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net972),
    .A1(net270),
    .A2(net1074),
    .A3(net831),
    .S0(net860),
    .S1(net973),
    .X(net273));
 sky130_fd_sc_hd__mux4_2 c467 (.A0(net162),
    .A1(net852),
    .A2(net2),
    .A3(clknet_1_1__leaf_net870),
    .S0(net522),
    .S1(net614),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net942),
    .A1(clknet_1_0__leaf_net253),
    .A2(net797),
    .A3(net1036),
    .S0(net905),
    .S1(net592),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(clknet_1_0__leaf_net133),
    .A1(net1049),
    .A2(clknet_1_1__leaf_net47),
    .A3(clknet_1_1__leaf_net898),
    .S0(net586),
    .S1(net649),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(clknet_1_1__leaf_net870),
    .A1(net96),
    .A2(net539),
    .A3(net905),
    .S0(net593),
    .S1(net640),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net809),
    .A1(net84),
    .A2(clknet_1_0__leaf_net115),
    .A3(net905),
    .S0(net593),
    .S1(net624),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net861),
    .A1(net942),
    .A2(net1000),
    .A3(net886),
    .S0(net1066),
    .S1(net652),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net841),
    .A1(net808),
    .A2(clknet_1_0__leaf_net893),
    .A3(net886),
    .S0(net614),
    .S1(net624),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net864),
    .A1(clknet_1_0__leaf_net112),
    .A2(clknet_1_0__leaf_net280),
    .A3(net1015),
    .S0(clknet_1_0__leaf_net899),
    .S1(net573),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_1__leaf_net280),
    .A1(clknet_1_1__leaf_net885),
    .A2(net948),
    .A3(net873),
    .S0(clknet_1_1__leaf_net898),
    .S1(net654),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(clknet_1_0__leaf_net115),
    .A1(net982),
    .A2(net640),
    .A3(net648),
    .S0(net650),
    .S1(net654),
    .X(net283));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net276),
    .A1(clknet_1_1__leaf_net59),
    .A2(net928),
    .A3(net1011),
    .S0(clknet_1_0__leaf_net902),
    .S1(net652),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net273),
    .A1(net1049),
    .A2(clknet_1_0__leaf_net62),
    .A3(net864),
    .S0(net949),
    .S1(net586),
    .X(net285));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net272),
    .A1(clknet_1_0__leaf_net280),
    .A2(clknet_1_0__leaf_net278),
    .A3(net844),
    .S0(net515),
    .S1(clknet_1_0__leaf_net890),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 c480 (.A0(net943),
    .A1(net854),
    .A2(net900),
    .A3(clknet_1_0__leaf_net280),
    .S0(clknet_1_0__leaf_net618),
    .S1(net655),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net1073),
    .A1(net951),
    .A2(clknet_1_0__leaf_net280),
    .A3(net854),
    .S0(clknet_1_0__leaf_net902),
    .S1(net656),
    .X(net895));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(net177),
    .A1(net283),
    .A2(net986),
    .A3(net900),
    .S0(net645),
    .S1(clknet_1_0__leaf_net657),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 c504 (.A0(net1014),
    .A1(net102),
    .A2(net1021),
    .A3(net1050),
    .S0(net980),
    .S1(net603),
    .X(net289));
 sky130_fd_sc_hd__mux4_2 c505 (.A0(net873),
    .A1(net1014),
    .A2(net992),
    .A3(net956),
    .S0(net289),
    .S1(net602),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 c506 (.A0(net1021),
    .A1(net955),
    .A2(net968),
    .A3(clknet_1_1__leaf_net544),
    .S0(net546),
    .S1(net604),
    .X(net291));
 sky130_fd_sc_hd__mux4_2 c507 (.A0(net951),
    .A1(net289),
    .A2(net290),
    .A3(net1017),
    .S0(net956),
    .S1(net962),
    .X(net292));
 sky130_fd_sc_hd__a41o_4 c508 (.A1(net998),
    .A2(net956),
    .A3(net503),
    .A4(net602),
    .B1(net605),
    .X(net293));
 sky130_fd_sc_hd__mux4_2 c509 (.A0(net1001),
    .A1(net1021),
    .A2(net293),
    .A3(net292),
    .S0(net992),
    .S1(net968),
    .X(net294));
 sky130_fd_sc_hd__a41o_1 c510 (.A1(net18),
    .A2(net945),
    .A3(net873),
    .A4(net293),
    .B1(clknet_1_0__leaf_net291),
    .X(net295));
 sky130_fd_sc_hd__mux4_1 c511 (.A0(net1021),
    .A1(net91),
    .A2(clknet_1_1__leaf_net291),
    .A3(net988),
    .S0(net294),
    .S1(net981),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c512 (.A0(net192),
    .A1(net871),
    .A2(clknet_1_1__leaf_net296),
    .A3(net956),
    .S0(net992),
    .S1(clknet_1_1__leaf_net291),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c513 (.A0(net91),
    .A1(net945),
    .A2(net290),
    .A3(clknet_1_1__leaf_net297),
    .S0(net601),
    .S1(net604),
    .X(net298));
 sky130_fd_sc_hd__a41o_1 c514 (.A1(net1014),
    .A2(clknet_1_1__leaf_net296),
    .A3(net110),
    .A4(clknet_1_1__leaf_net297),
    .B1(net289),
    .X(net299));
 sky130_fd_sc_hd__sdfbbn_1 c515 (.CLK_N(clknet_leaf_18_clk),
    .D(clknet_1_0__leaf_net296),
    .RESET_B(net293),
    .SCD(clknet_1_1__leaf_net299),
    .SCE(clknet_1_1__leaf_net297),
    .SET_B(clknet_1_1__leaf_net204),
    .Q(net301),
    .Q_N(net300));
 sky130_fd_sc_hd__mux4_1 c516 (.A0(net301),
    .A1(clknet_1_1__leaf_net299),
    .A2(net945),
    .A3(net289),
    .S0(net1008),
    .S1(clknet_1_1__leaf_net291),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net289),
    .A1(net293),
    .A2(net777),
    .A3(clknet_1_1__leaf_net291),
    .S0(clknet_1_1__leaf_net299),
    .S1(net660),
    .X(net303));
 sky130_fd_sc_hd__mux4_1 c518 (.A0(net290),
    .A1(net189),
    .A2(net300),
    .A3(clknet_1_1__leaf_net299),
    .S0(net871),
    .S1(net1039),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net196),
    .A1(net192),
    .A2(clknet_1_1__leaf_net296),
    .A3(net300),
    .S0(clknet_1_1__leaf_net299),
    .S1(net1017),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c520 (.A0(clknet_1_1__leaf_net299),
    .A1(clknet_1_1__leaf_net295),
    .A2(clknet_1_0__leaf_net296),
    .A3(net981),
    .S0(clknet_1_1__leaf_net596),
    .S1(net664),
    .X(net306));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(net301),
    .A1(net91),
    .A2(net661),
    .A3(net663),
    .S0(net664),
    .S1(net665),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net307),
    .A1(net873),
    .A2(net825),
    .A3(net662),
    .S0(net664),
    .S1(net665),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 c523 (.A0(net307),
    .A1(net292),
    .A2(net290),
    .A3(net503),
    .S0(net661),
    .S1(net665),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net1012),
    .A1(clknet_1_1__leaf_net291),
    .A2(net308),
    .A3(net307),
    .S0(net664),
    .S1(net665),
    .X(net310));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(clknet_1_1__leaf_net295),
    .A1(net294),
    .A2(net1052),
    .A3(clknet_1_1__leaf_net114),
    .S0(net525),
    .S1(clknet_1_1__leaf_net616),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net208),
    .A1(clknet_1_0__leaf_net204),
    .A2(net289),
    .A3(clknet_1_0__leaf_net291),
    .S0(net960),
    .S1(net993),
    .X(net312));
 sky130_fd_sc_hd__mux4_1 c527 (.A0(net953),
    .A1(net1006),
    .A2(net998),
    .A3(net525),
    .S0(clknet_1_0__leaf_net617),
    .S1(net619),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c528 (.A0(net191),
    .A1(net6),
    .A2(net953),
    .A3(net799),
    .S0(net525),
    .S1(net620),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 c529 (.A0(clknet_1_0__leaf_net296),
    .A1(clknet_1_0__leaf_net313),
    .A2(net802),
    .A3(clknet_1_1__leaf_net883),
    .S0(net915),
    .S1(net869),
    .X(net315));
 sky130_fd_sc_hd__mux4_1 c530 (.A0(net33),
    .A1(clknet_1_1__leaf_net299),
    .A2(clknet_1_0__leaf_net297),
    .A3(net1070),
    .S0(net525),
    .S1(net666),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c531 (.A0(clknet_1_0__leaf_net313),
    .A1(net994),
    .A2(clknet_1_0__leaf_net299),
    .A3(net993),
    .S0(net956),
    .S1(clknet_1_1__leaf_net617),
    .X(net317));
 sky130_fd_sc_hd__mux4_1 c532 (.A0(net314),
    .A1(net915),
    .A2(clknet_1_0__leaf_net207),
    .A3(clknet_1_0__leaf_net297),
    .S0(net992),
    .S1(net561),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c533 (.A0(clknet_1_1__leaf_net222),
    .A1(net1050),
    .A2(net802),
    .A3(net981),
    .S0(net668),
    .S1(net672),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 c534 (.A0(net293),
    .A1(net18),
    .A2(net33),
    .A3(net608),
    .S0(clknet_1_0__leaf_net617),
    .S1(net672),
    .X(net320));
 sky130_fd_sc_hd__mux4_2 c535 (.A0(net1031),
    .A1(net994),
    .A2(net552),
    .A3(net620),
    .S0(net667),
    .S1(net673),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c536 (.A0(net945),
    .A1(net300),
    .A2(net666),
    .A3(net667),
    .S0(net670),
    .S1(net673),
    .X(net322));
 sky130_fd_sc_hd__mux4_1 c537 (.A0(net322),
    .A1(clknet_1_1__leaf_net312),
    .A2(net292),
    .A3(net956),
    .S0(net873),
    .S1(net110),
    .X(net323));
 sky130_fd_sc_hd__mux4_1 c538 (.A0(net789),
    .A1(net1052),
    .A2(net189),
    .A3(net960),
    .S0(net599),
    .S1(clknet_1_0__leaf_net675),
    .X(net324));
 sky130_fd_sc_hd__mux4_1 c539 (.A0(clknet_1_0__leaf_net324),
    .A1(net322),
    .A2(net33),
    .A3(net1001),
    .S0(net667),
    .S1(clknet_1_0__leaf_net675),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c540 (.A0(clknet_1_0__leaf_net297),
    .A1(clknet_1_1__leaf_net324),
    .A2(net803),
    .A3(clknet_1_1__leaf_net883),
    .S0(net554),
    .S1(clknet_1_1__leaf_net888),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c541 (.A0(net294),
    .A1(clknet_1_1__leaf_net883),
    .A2(net608),
    .A3(net673),
    .S0(clknet_1_1__leaf_net888),
    .S1(clknet_1_0__leaf_net676),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 c542 (.A0(net321),
    .A1(clknet_1_0__leaf_net324),
    .A2(clknet_1_0__leaf_net299),
    .A3(clknet_1_0__leaf_net313),
    .S0(clknet_1_1__leaf_net675),
    .S1(clknet_1_0__leaf_net676),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 c543 (.A0(net506),
    .A1(clknet_1_1__leaf_net544),
    .A2(clknet_1_1__leaf_net596),
    .A3(net672),
    .S0(net673),
    .S1(net674),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c544 (.A0(clknet_1_1__leaf_net329),
    .A1(net322),
    .A2(clknet_1_1__leaf_net562),
    .A3(net666),
    .S0(clknet_1_1__leaf_net888),
    .S1(net678),
    .X(net330));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(clknet_1_0__leaf_net329),
    .A1(net506),
    .A2(net673),
    .A3(net674),
    .S0(clknet_1_0__leaf_net676),
    .S1(net677),
    .X(net331));
 sky130_fd_sc_hd__sdfbbn_1 c546 (.CLK_N(clknet_leaf_34_clk),
    .D(clknet_1_0__leaf_net299),
    .RESET_B(clknet_1_0__leaf_net295),
    .SCD(clknet_1_0__leaf_net883),
    .SCE(net510),
    .SET_B(net674),
    .Q(net333),
    .Q_N(net332));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(clknet_1_0__leaf_net312),
    .A1(net18),
    .A2(net994),
    .A3(net1038),
    .S0(net564),
    .S1(net569),
    .X(net334));
 sky130_fd_sc_hd__mux4_2 c548 (.A0(net791),
    .A1(net1009),
    .A2(net782),
    .A3(net556),
    .S0(net631),
    .S1(net669),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(clknet_1_0__leaf_net234),
    .A1(net790),
    .A2(net1027),
    .A3(net772),
    .S0(net612),
    .S1(net673),
    .X(net336));
 sky130_fd_sc_hd__mux4_1 c550 (.A0(clknet_1_1__leaf_net229),
    .A1(net984),
    .A2(net557),
    .A3(net565),
    .S0(net569),
    .S1(net680),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c551 (.A0(clknet_1_0__leaf_net324),
    .A1(clknet_1_1__leaf_net295),
    .A2(net1017),
    .A3(net1100),
    .S0(net572),
    .S1(net681),
    .X(net338));
 sky130_fd_sc_hd__mux4_1 c552 (.A0(net333),
    .A1(clknet_1_0__leaf_net331),
    .A2(net18),
    .A3(net569),
    .S0(net572),
    .S1(net665),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c553 (.A0(clknet_1_0__leaf_net204),
    .A1(net239),
    .A2(net1007),
    .A3(net564),
    .S0(net572),
    .S1(net681),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c554 (.A0(net945),
    .A1(clknet_1_1__leaf_net233),
    .A2(clknet_1_0__leaf_net247),
    .A3(clknet_1_0__leaf_net204),
    .S0(net321),
    .S1(net1014),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c555 (.A0(net301),
    .A1(net321),
    .A2(clknet_1_1__leaf_net337),
    .A3(net510),
    .S0(net564),
    .S1(net572),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c556 (.A0(clknet_1_0__leaf_net331),
    .A1(clknet_1_0__leaf_net312),
    .A2(clknet_1_0__leaf_net299),
    .A3(net632),
    .S0(net673),
    .S1(net684),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 c557 (.A0(clknet_1_0__leaf_net234),
    .A1(clknet_1_1__leaf_net339),
    .A2(net518),
    .A3(net564),
    .S0(net682),
    .S1(net685),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 c558 (.A0(net962),
    .A1(net39),
    .A2(net818),
    .A3(net607),
    .S0(net681),
    .S1(net686),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 c559 (.A0(clknet_1_0__leaf_net331),
    .A1(net345),
    .A2(net1070),
    .A3(net292),
    .S0(net610),
    .S1(net686),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(clknet_1_0__leaf_net346),
    .A1(clknet_1_0__leaf_net340),
    .A2(clknet_1_0__leaf_net299),
    .A3(clknet_1_0__leaf_net544),
    .S0(net565),
    .S1(net685),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 c561 (.A0(clknet_1_0__leaf_net339),
    .A1(net1000),
    .A2(net915),
    .A3(net982),
    .S0(net554),
    .S1(net687),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 c562 (.A0(net321),
    .A1(net345),
    .A2(clknet_1_0__leaf_net346),
    .A3(net605),
    .S0(net686),
    .S1(net687),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(clknet_1_0__leaf_net337),
    .A1(net1003),
    .A2(net957),
    .A3(net871),
    .S0(net632),
    .S1(net683),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c564 (.A0(net350),
    .A1(net345),
    .A2(clknet_1_1__leaf_net348),
    .A3(net321),
    .S0(net988),
    .S1(net1014),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net345),
    .A1(clknet_1_0__leaf_net324),
    .A2(clknet_1_1__leaf_net346),
    .A3(clknet_1_1__leaf_net331),
    .S0(clknet_1_0__leaf_net298),
    .S1(net816),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(clknet_1_1__leaf_net340),
    .A1(clknet_1_1__leaf_net247),
    .A2(net40),
    .A3(net777),
    .S0(net669),
    .S1(net687),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c567 (.A0(clknet_1_0__leaf_net233),
    .A1(net928),
    .A2(clknet_1_0__leaf_net295),
    .A3(net506),
    .S0(net605),
    .S1(net692),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net790),
    .A1(net957),
    .A2(net532),
    .A3(clknet_1_1__leaf_net638),
    .S0(net682),
    .S1(net687),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c569 (.A0(net826),
    .A1(net994),
    .A2(clknet_1_0__leaf_net883),
    .A3(net1053),
    .S0(clknet_1_0__leaf_net544),
    .S1(clknet_1_0__leaf_net638),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net355),
    .A1(net333),
    .A2(clknet_1_0__leaf_net291),
    .A3(net988),
    .S0(net844),
    .S1(clknet_1_1__leaf_net638),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c571 (.A0(net787),
    .A1(net1028),
    .A2(clknet_1_1__leaf_net47),
    .A3(net645),
    .S0(net678),
    .S1(net685),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c572 (.A0(net790),
    .A1(net113),
    .A2(net531),
    .A3(net573),
    .S0(net677),
    .S1(net695),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(clknet_1_0__leaf_net226),
    .A1(clknet_1_1__leaf_net257),
    .A2(net518),
    .A3(net521),
    .S0(net605),
    .S1(clknet_1_0__leaf_net696),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c574 (.A0(clknet_1_0__leaf_net295),
    .A1(net110),
    .A2(net844),
    .A3(clknet_1_1__leaf_net165),
    .S0(net631),
    .S1(net688),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(clknet_1_0__leaf_net220),
    .A1(clknet_1_0__leaf_net243),
    .A2(clknet_1_0__leaf_net342),
    .A3(clknet_1_0__leaf_net544),
    .S0(net614),
    .S1(clknet_1_0__leaf_net696),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net819),
    .A1(net1001),
    .A2(clknet_1_1__leaf_net47),
    .A3(clknet_1_0__leaf_net544),
    .S0(net646),
    .S1(net694),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(clknet_1_0__leaf_net363),
    .A1(clknet_1_0__leaf_net220),
    .A2(net1078),
    .A3(net787),
    .S0(clknet_1_0__leaf_net158),
    .S1(net687),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(clknet_1_0__leaf_net220),
    .A1(net801),
    .A2(net1051),
    .A3(clknet_1_1__leaf_net363),
    .S0(net682),
    .S1(net698),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net986),
    .A1(net332),
    .A2(clknet_1_0__leaf_net291),
    .A3(net636),
    .S0(net679),
    .S1(net702),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net831),
    .A1(clknet_1_0__leaf_net882),
    .A2(net527),
    .A3(net532),
    .S0(clknet_1_1__leaf_net581),
    .S1(clknet_1_1__leaf_net696),
    .X(net877));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(clknet_1_1__leaf_net357),
    .A1(net951),
    .A2(net518),
    .A3(net537),
    .S0(clknet_1_0__leaf_net888),
    .S1(net701),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(clknet_1_1__leaf_net357),
    .A1(net791),
    .A2(net799),
    .A3(clknet_1_0__leaf_net544),
    .S0(clknet_1_1__leaf_net696),
    .S1(net700),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net52),
    .A1(net1075),
    .A2(net844),
    .A3(clknet_1_0__leaf_net367),
    .S0(clknet_1_0__leaf_net348),
    .S1(net946),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net988),
    .A1(net957),
    .A2(clknet_1_0__leaf_net357),
    .A3(clknet_1_1__leaf_net257),
    .S0(net52),
    .S1(net697),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(clknet_1_0__leaf_net357),
    .A1(clknet_1_0__leaf_net368),
    .A2(net527),
    .A3(net569),
    .S0(net625),
    .S1(net703),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(clknet_1_1__leaf_net367),
    .A1(net827),
    .A2(net819),
    .A3(clknet_1_0__leaf_net363),
    .S0(net986),
    .S1(net973),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_1__leaf_net158),
    .A1(net1079),
    .A2(net1035),
    .A3(clknet_1_1__leaf_net372),
    .S0(clknet_1_0__leaf_net368),
    .S1(net986),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net1051),
    .A1(clknet_1_0__leaf_net342),
    .A2(net2),
    .A3(net844),
    .S0(net947),
    .S1(net647),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net1019),
    .A1(net799),
    .A2(net1015),
    .A3(clknet_1_0__leaf_net883),
    .S0(net791),
    .S1(net861),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net848),
    .A1(clknet_1_0__leaf_net282),
    .A2(net1074),
    .A3(clknet_1_1__leaf_net178),
    .S0(net802),
    .S1(net679),
    .X(net376));
 sky130_fd_sc_hd__mux4_2 c591 (.A0(net808),
    .A1(net802),
    .A2(net1051),
    .A3(net1008),
    .S0(net872),
    .S1(net705),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net827),
    .A1(net831),
    .A2(net377),
    .A3(clknet_1_1__leaf_net178),
    .S0(net589),
    .S1(net647),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net369),
    .A1(net1074),
    .A2(clknet_1_0__leaf_net883),
    .A3(clknet_1_1__leaf_net282),
    .S0(net995),
    .S1(net957),
    .X(net379));
 sky130_fd_sc_hd__mux4_2 c594 (.A0(net873),
    .A1(net973),
    .A2(net951),
    .A3(net658),
    .S0(net680),
    .S1(net699),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(clknet_1_1__leaf_net78),
    .A1(clknet_1_1__leaf_net278),
    .A2(net380),
    .A3(net827),
    .S0(net947),
    .S1(net871),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net866),
    .A1(net949),
    .A2(net583),
    .A3(net588),
    .S0(net645),
    .S1(net693),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net866),
    .A1(net366),
    .A2(net860),
    .A3(clknet_1_1__leaf_net165),
    .S0(net645),
    .S1(net659),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net380),
    .A1(net1015),
    .A2(net1019),
    .A3(clknet_1_0__leaf_net883),
    .S0(net522),
    .S1(net706),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 c599 (.A0(net861),
    .A1(net957),
    .A2(net1000),
    .A3(net582),
    .S0(net659),
    .S1(net706),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(clknet_1_1__leaf_net47),
    .A1(net1004),
    .A2(net377),
    .A3(net565),
    .S0(net583),
    .S1(net709),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net371),
    .A1(net944),
    .A2(net871),
    .A3(net1075),
    .S0(clknet_1_0__leaf_net657),
    .S1(net705),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net2),
    .A1(net790),
    .A2(net802),
    .A3(net1000),
    .S0(net878),
    .S1(clknet_1_0__leaf_net618),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net1000),
    .A1(clknet_1_0__leaf_net243),
    .A2(clknet_1_0__leaf_net388),
    .A3(net600),
    .S0(net614),
    .S1(net710),
    .X(net389));
 sky130_fd_sc_hd__mux4_2 c604 (.A0(net380),
    .A1(net944),
    .A2(net573),
    .A3(net701),
    .S0(net710),
    .S1(net711),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(clknet_1_0__leaf_net348),
    .A1(clknet_1_1__leaf_net388),
    .A2(net866),
    .A3(net645),
    .S0(clknet_1_1__leaf_net657),
    .S1(net678),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(clknet_1_0__leaf_net388),
    .A1(clknet_1_0__leaf_net882),
    .A2(net377),
    .A3(net1014),
    .S0(net710),
    .S1(net711),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(clknet_1_1__leaf_net165),
    .A1(net382),
    .A2(net392),
    .A3(clknet_1_1__leaf_net178),
    .S0(net1074),
    .S1(net653),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(clknet_1_1__leaf_net178),
    .A1(clknet_1_0__leaf_net883),
    .A2(net514),
    .A3(net639),
    .S0(net706),
    .S1(net712),
    .X(net394));
 sky130_fd_sc_hd__mux4_2 c630 (.A0(net309),
    .A1(net962),
    .A2(net187),
    .A3(net308),
    .S0(net980),
    .S1(net599),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net308),
    .A1(net956),
    .A2(net309),
    .A3(clknet_1_1__leaf_net310),
    .S0(net777),
    .S1(net503),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(clknet_1_0__leaf_net310),
    .A1(net39),
    .A2(net999),
    .A3(net992),
    .S0(net309),
    .S1(net503),
    .X(net397));
 sky130_fd_sc_hd__mux4_2 c633 (.A0(net7),
    .A1(net953),
    .A2(net962),
    .A3(net988),
    .S0(net1017),
    .S1(net395),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(clknet_1_1__leaf_net396),
    .A1(clknet_1_1__leaf_net204),
    .A2(net995),
    .A3(clknet_1_1__leaf_net291),
    .S0(net992),
    .S1(net663),
    .X(net399));
 sky130_fd_sc_hd__mux4_1 c635 (.A0(net951),
    .A1(net1048),
    .A2(clknet_1_0__leaf_net399),
    .A3(net189),
    .S0(net398),
    .S1(net992),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net190),
    .A1(net189),
    .A2(clknet_1_1__leaf_net399),
    .A3(net984),
    .S0(net995),
    .S1(clknet_1_1__leaf_net598),
    .X(net401));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net398),
    .A1(net293),
    .A2(net993),
    .A3(net956),
    .S0(net1001),
    .S1(net714),
    .X(net402));
 sky130_fd_sc_hd__mux4_1 c638 (.A0(net953),
    .A1(net1001),
    .A2(clknet_1_1__leaf_net399),
    .A3(net1015),
    .S0(net503),
    .S1(net981),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 c639 (.A0(net188),
    .A1(net102),
    .A2(clknet_1_1__leaf_net299),
    .A3(net999),
    .S0(net981),
    .S1(net599),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 c640 (.A0(net993),
    .A1(clknet_1_0__leaf_net310),
    .A2(clknet_1_1__leaf_net397),
    .A3(net973),
    .S0(net545),
    .S1(net719),
    .X(net405));
 sky130_fd_sc_hd__mux4_1 c641 (.A0(clknet_1_1__leaf_net299),
    .A1(net402),
    .A2(clknet_1_1__leaf_net396),
    .A3(clknet_1_1__leaf_net405),
    .S0(clknet_1_1__leaf_net598),
    .S1(net716),
    .X(net406));
 sky130_fd_sc_hd__mux4_1 c642 (.A0(net402),
    .A1(net988),
    .A2(clknet_1_1__leaf_net310),
    .A3(net960),
    .S0(net398),
    .S1(net499),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 c643 (.A0(clknet_1_1__leaf_net396),
    .A1(net293),
    .A2(net294),
    .A3(net395),
    .S0(net499),
    .S1(net720),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(clknet_1_1__leaf_net397),
    .A1(net309),
    .A2(net546),
    .A3(net716),
    .S0(net718),
    .S1(net721),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 c645 (.A0(clknet_1_1__leaf_net408),
    .A1(net402),
    .A2(net1001),
    .A3(clknet_1_1__leaf_net399),
    .S0(net953),
    .S1(net721),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 c646 (.A0(clknet_1_1__leaf_net409),
    .A1(clknet_1_1__leaf_net204),
    .A2(net956),
    .A3(clknet_1_0__leaf_net408),
    .S0(net720),
    .S1(net722),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c647 (.A0(net402),
    .A1(net190),
    .A2(net7),
    .A3(net500),
    .S0(net599),
    .S1(net721),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 c648 (.A0(clknet_1_1__leaf_net399),
    .A1(clknet_1_0__leaf_net408),
    .A2(clknet_1_0__leaf_net409),
    .A3(net503),
    .S0(net721),
    .S1(net723),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(clknet_1_1__leaf_net411),
    .A1(clknet_1_1__leaf_net396),
    .A2(net102),
    .A3(net720),
    .S0(net721),
    .S1(net723),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(net963),
    .A1(clknet_1_0__leaf_net409),
    .A2(clknet_1_1__leaf_net397),
    .A3(net500),
    .S0(net722),
    .S1(net724),
    .X(net415));
 sky130_fd_sc_hd__mux4_1 c651 (.A0(net188),
    .A1(clknet_1_1__leaf_net405),
    .A2(clknet_1_1__leaf_net331),
    .A3(net294),
    .S0(net984),
    .S1(net615),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c652 (.A0(clknet_1_1__leaf_net204),
    .A1(clknet_1_1__leaf_net405),
    .A2(clknet_1_0__leaf_net397),
    .A3(net973),
    .S0(net1070),
    .S1(clknet_1_1__leaf_net676),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c653 (.A0(net787),
    .A1(net395),
    .A2(clknet_1_1__leaf_net204),
    .A3(net6),
    .S0(clknet_1_1__leaf_net888),
    .S1(net723),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 c654 (.A0(net395),
    .A1(net314),
    .A2(net781),
    .A3(net521),
    .S0(net608),
    .S1(net869),
    .X(net419));
 sky130_fd_sc_hd__mux4_1 c655 (.A0(clknet_1_0__leaf_net415),
    .A1(net292),
    .A2(net988),
    .A3(net561),
    .S0(clknet_1_1__leaf_net596),
    .S1(net715),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c656 (.A0(net782),
    .A1(net314),
    .A2(clknet_1_1__leaf_net888),
    .A3(clknet_1_1__leaf_net676),
    .S0(net723),
    .S1(net724),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(clknet_1_0__leaf_net397),
    .A1(net787),
    .A2(net187),
    .A3(net1039),
    .S0(net609),
    .S1(net718),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(clknet_1_0__leaf_net397),
    .A1(clknet_1_0__leaf_net418),
    .A2(net101),
    .A3(net39),
    .S0(net664),
    .S1(net726),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net802),
    .A1(net110),
    .A2(clknet_1_0__leaf_net415),
    .A3(net995),
    .S0(net552),
    .S1(net609),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 c660 (.A0(clknet_1_1__leaf_net417),
    .A1(clknet_1_1__leaf_net207),
    .A2(clknet_1_1__leaf_net298),
    .A3(net995),
    .S0(net714),
    .S1(net717),
    .X(net425));
 sky130_fd_sc_hd__mux4_1 c661 (.A0(clknet_1_1__leaf_net298),
    .A1(net801),
    .A2(clknet_1_1__leaf_net226),
    .A3(clknet_1_1__leaf_net405),
    .S0(net724),
    .S1(net729),
    .X(net426));
 sky130_fd_sc_hd__mux4_1 c662 (.A0(net218),
    .A1(net289),
    .A2(net993),
    .A3(net801),
    .S0(net521),
    .S1(net730),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c663 (.A0(net189),
    .A1(net947),
    .A2(clknet_1_0__leaf_net396),
    .A3(net989),
    .S0(net505),
    .S1(clknet_1_1__leaf_net888),
    .X(net428));
 sky130_fd_sc_hd__mux4_1 c664 (.A0(net294),
    .A1(net977),
    .A2(clknet_1_1__leaf_net207),
    .A3(net963),
    .S0(net730),
    .S1(net731),
    .X(net429));
 sky130_fd_sc_hd__mux4_1 c665 (.A0(clknet_1_1__leaf_net396),
    .A1(clknet_1_1__leaf_net428),
    .A2(net505),
    .A3(net719),
    .S0(net723),
    .S1(net725),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 c666 (.A0(net802),
    .A1(clknet_1_0__leaf_net429),
    .A2(net427),
    .A3(net521),
    .S0(net552),
    .S1(net729),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 c667 (.A0(clknet_1_1__leaf_net428),
    .A1(net715),
    .A2(net726),
    .A3(net728),
    .S0(net729),
    .S1(net731),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c668 (.A0(clknet_1_1__leaf_net418),
    .A1(clknet_1_1__leaf_net207),
    .A2(net993),
    .A3(clknet_1_1__leaf_net226),
    .S0(clknet_1_0__leaf_net428),
    .S1(clknet_1_1__leaf_net733),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 c669 (.A0(clknet_1_0__leaf_net399),
    .A1(net427),
    .A2(clknet_1_1__leaf_net429),
    .A3(net505),
    .S0(clknet_1_1__leaf_net596),
    .S1(clknet_1_0__leaf_net733),
    .X(net434));
 sky130_fd_sc_hd__mux4_1 c670 (.A0(clknet_1_0__leaf_net428),
    .A1(net427),
    .A2(clknet_1_0__leaf_net417),
    .A3(net110),
    .S0(net729),
    .S1(net737),
    .X(net435));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(clknet_1_1__leaf_net415),
    .A1(net289),
    .A2(net723),
    .A3(net727),
    .S0(net737),
    .S1(net739),
    .X(net436));
 sky130_fd_sc_hd__mux4_1 c672 (.A0(net993),
    .A1(net947),
    .A2(net1001),
    .A3(net187),
    .S0(clknet_1_1__leaf_net416),
    .S1(clknet_1_1__leaf_net734),
    .X(net437));
 sky130_fd_sc_hd__mux4_1 c673 (.A0(clknet_1_1__leaf_net411),
    .A1(net335),
    .A2(net572),
    .A3(net731),
    .S0(net736),
    .S1(net740),
    .X(net438));
 sky130_fd_sc_hd__mux4_1 c674 (.A0(clknet_1_1__leaf_net114),
    .A1(net110),
    .A2(net973),
    .A3(net671),
    .S0(net717),
    .S1(net741),
    .X(net439));
 sky130_fd_sc_hd__mux4_1 c675 (.A0(net43),
    .A1(net239),
    .A2(net995),
    .A3(net674),
    .S0(clknet_1_0__leaf_net734),
    .S1(net743),
    .X(net440));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net293),
    .A1(net1007),
    .A2(net505),
    .A3(net626),
    .S0(net689),
    .S1(net735),
    .X(net441));
 sky130_fd_sc_hd__mux4_1 c677 (.A0(net289),
    .A1(clknet_1_0__leaf_net396),
    .A2(net607),
    .A3(clknet_1_1__leaf_net888),
    .S0(net730),
    .S1(net737),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net102),
    .A1(net1101),
    .A2(net43),
    .A3(clknet_1_1__leaf_net442),
    .S0(net977),
    .S1(net730),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net791),
    .A1(net1007),
    .A2(net1012),
    .A3(net626),
    .S0(clknet_1_0__leaf_net888),
    .S1(net722),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(clknet_1_1__leaf_net234),
    .A1(clknet_1_0__leaf_net396),
    .A2(clknet_1_0__leaf_net299),
    .A3(net691),
    .S0(net692),
    .S1(net722),
    .X(net445));
 sky130_fd_sc_hd__mux4_1 c681 (.A0(clknet_1_1__leaf_net241),
    .A1(clknet_1_1__leaf_net442),
    .A2(net1017),
    .A3(clknet_1_0__leaf_net204),
    .S0(net722),
    .S1(clknet_1_0__leaf_net732),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c682 (.A0(clknet_1_0__leaf_net399),
    .A1(net963),
    .A2(clknet_1_0__leaf_net204),
    .A3(clknet_1_0__leaf_net396),
    .S0(net773),
    .S1(clknet_1_0__leaf_net888),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c683 (.A0(net443),
    .A1(clknet_1_1__leaf_net446),
    .A2(clknet_1_1__leaf_net142),
    .A3(clknet_1_0__leaf_net396),
    .S0(clknet_1_1__leaf_net562),
    .S1(net716),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net26),
    .A1(net773),
    .A2(net572),
    .A3(net717),
    .S0(clknet_1_1__leaf_net732),
    .S1(net745),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c685 (.A0(net26),
    .A1(net335),
    .A2(net504),
    .A3(clknet_1_0__leaf_net888),
    .S0(net738),
    .S1(net744),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(clknet_1_0__leaf_net298),
    .A1(clknet_1_1__leaf_net313),
    .A2(net335),
    .A3(net818),
    .S0(net774),
    .S1(net599),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c687 (.A0(net449),
    .A1(net230),
    .A2(clknet_1_1__leaf_net142),
    .A3(net968),
    .S0(clknet_1_1__leaf_net562),
    .S1(net572),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c688 (.A0(clknet_1_1__leaf_net142),
    .A1(net1007),
    .A2(clknet_1_1__leaf_net452),
    .A3(net504),
    .S0(net508),
    .S1(net674),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net453),
    .A1(clknet_1_1__leaf_net452),
    .A2(net26),
    .A3(net670),
    .S0(net722),
    .S1(net744),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c690 (.A0(net292),
    .A1(clknet_1_1__leaf_net313),
    .A2(clknet_1_0__leaf_net399),
    .A3(clknet_1_1__leaf_net452),
    .S0(clknet_1_1__leaf_net442),
    .S1(net993),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c691 (.A0(net454),
    .A1(net335),
    .A2(clknet_1_1__leaf_net452),
    .A3(net690),
    .S0(net730),
    .S1(net742),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(clknet_1_0__leaf_net452),
    .A1(net1004),
    .A2(net665),
    .A3(net671),
    .S0(net691),
    .S1(net748),
    .X(net457));
 sky130_fd_sc_hd__mux4_1 c693 (.A0(net40),
    .A1(net963),
    .A2(net1008),
    .A3(clknet_1_1__leaf_net226),
    .S0(clknet_1_0__leaf_net405),
    .S1(clknet_1_0__leaf_net442),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c694 (.A0(clknet_1_1__leaf_net207),
    .A1(net439),
    .A2(clknet_1_1__leaf_net342),
    .A3(net600),
    .S0(net633),
    .S1(net738),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c695 (.A0(net1008),
    .A1(clknet_1_0__leaf_net452),
    .A2(clknet_1_1__leaf_net349),
    .A3(net625),
    .S0(net644),
    .S1(net731),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net113),
    .A1(net1047),
    .A2(net1004),
    .A3(net787),
    .S0(net646),
    .S1(clknet_1_0__leaf_net888),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c697 (.A0(clknet_1_0__leaf_net446),
    .A1(net441),
    .A2(net1040),
    .A3(net187),
    .S0(net704),
    .S1(net741),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 c698 (.A0(net441),
    .A1(net831),
    .A2(net1036),
    .A3(net522),
    .S0(net633),
    .S1(net869),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c699 (.A0(clknet_1_0__leaf_net405),
    .A1(clknet_1_1__leaf_net368),
    .A2(net982),
    .A3(net552),
    .S0(net646),
    .S1(net744),
    .X(net464));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(clknet_1_0__leaf_net291),
    .A1(net239),
    .A2(net293),
    .A3(clknet_1_0__leaf_net142),
    .S0(net645),
    .S1(net721),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(clknet_1_1__leaf_net226),
    .A1(clknet_1_1__leaf_net142),
    .A2(clknet_1_1__leaf_net444),
    .A3(net558),
    .S0(net747),
    .S1(clknet_1_1__leaf_net752),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c702 (.A0(clknet_1_0__leaf_net405),
    .A1(net40),
    .A2(net1015),
    .A3(net671),
    .S0(net750),
    .S1(clknet_1_1__leaf_net754),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(clknet_1_1__leaf_net467),
    .A1(net110),
    .A2(net464),
    .A3(net463),
    .S0(net188),
    .S1(clknet_1_1__leaf_net753),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net1040),
    .A1(net963),
    .A2(net1008),
    .A3(clknet_1_1__leaf_net62),
    .S0(net633),
    .S1(net743),
    .X(net469));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(clknet_1_0__leaf_net416),
    .A1(clknet_1_1__leaf_net422),
    .A2(net40),
    .A3(net818),
    .S0(clknet_1_0__leaf_net442),
    .S1(net463),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net988),
    .A1(clknet_1_0__leaf_net405),
    .A2(net689),
    .A3(net703),
    .S0(net729),
    .S1(net741),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(clknet_1_1__leaf_net368),
    .A1(net110),
    .A2(clknet_1_0__leaf_net422),
    .A3(clknet_1_1__leaf_net581),
    .S0(net688),
    .S1(net703),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net110),
    .A1(net643),
    .A2(net689),
    .A3(net692),
    .S0(net721),
    .S1(net738),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net463),
    .A1(net1004),
    .A2(clknet_1_0__leaf_net452),
    .A3(net579),
    .S0(net729),
    .S1(net748),
    .X(net474));
 sky130_fd_sc_hd__mux4_1 c710 (.A0(net473),
    .A1(net984),
    .A2(clknet_1_1__leaf_net226),
    .A3(clknet_1_0__leaf_net467),
    .S0(clknet_1_0__leaf_net416),
    .S1(net565),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net818),
    .A1(net474),
    .A2(net839),
    .A3(clknet_1_1__leaf_net207),
    .S0(net982),
    .S1(net744),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(clknet_1_1__leaf_net476),
    .A1(net645),
    .A2(net692),
    .A3(net731),
    .S0(net751),
    .S1(net759),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(net801),
    .A1(clknet_1_0__leaf_net476),
    .A2(net839),
    .A3(net984),
    .S0(net721),
    .S1(net760),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net440),
    .A1(clknet_1_0__leaf_net411),
    .A2(net472),
    .A3(net386),
    .S0(net561),
    .S1(net692),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net184),
    .A1(net378),
    .A2(net522),
    .A3(net982),
    .S0(net625),
    .S1(net694),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(clknet_1_0__leaf_net299),
    .A1(net1036),
    .A2(net1001),
    .A3(clknet_1_1__leaf_net62),
    .S0(net561),
    .S1(net759),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net995),
    .A1(net799),
    .A2(net831),
    .A3(net583),
    .S0(net692),
    .S1(net705),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net1075),
    .A1(net457),
    .A2(net391),
    .A3(clknet_1_0__leaf_net349),
    .S0(net645),
    .S1(clknet_1_0__leaf_net752),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(net1036),
    .A1(net1007),
    .A2(net501),
    .A3(net579),
    .S0(clknet_1_1__leaf_net657),
    .S1(net749),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_0__leaf_net446),
    .A1(clknet_1_0__leaf_net444),
    .A2(net951),
    .A3(net565),
    .S0(clknet_1_0__leaf_net754),
    .S1(net763),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(clknet_1_1__leaf_net62),
    .A1(net1019),
    .A2(net860),
    .A3(net774),
    .S0(net713),
    .S1(net762),
    .X(net486));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net951),
    .A1(clknet_1_1__leaf_net142),
    .A2(net377),
    .A3(net484),
    .S0(net640),
    .S1(net763),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(clknet_1_0__leaf_net442),
    .A1(net839),
    .A2(net858),
    .A3(net565),
    .S0(net595),
    .S1(net758),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(clknet_1_1__leaf_net342),
    .A1(net1053),
    .A2(net860),
    .A3(net982),
    .S0(net579),
    .S1(net756),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net1004),
    .A1(net465),
    .A2(net385),
    .A3(net1014),
    .S0(net982),
    .S1(net640),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net487),
    .A1(net947),
    .A2(net450),
    .A3(net488),
    .S0(clknet_1_1__leaf_net62),
    .S1(net766),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net844),
    .A1(net482),
    .A2(net879),
    .A3(net653),
    .S0(net764),
    .S1(net767),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net973),
    .A1(net839),
    .A2(net502),
    .A3(net982),
    .S0(net561),
    .S1(net600),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_0__leaf_net372),
    .A1(clknet_1_0__leaf_net349),
    .A2(net1075),
    .A3(net492),
    .S0(clknet_1_0__leaf_net411),
    .S1(net711),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net831),
    .A1(net1053),
    .A2(net490),
    .A3(net694),
    .S0(net761),
    .S1(net769),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net858),
    .A1(net1012),
    .A2(net746),
    .A3(clknet_1_0__leaf_net753),
    .S0(net755),
    .S1(net768),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net791),
    .A1(net774),
    .A2(net471),
    .A3(net495),
    .S0(net707),
    .S1(net708),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net230),
    .A1(net973),
    .A2(net493),
    .A3(net463),
    .S0(net496),
    .S1(net742),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(net1007),
    .A1(net498),
    .A2(net745),
    .A3(net757),
    .S0(net765),
    .S1(net770));
 sky130_fd_sc_hd__dfrbp_1 merge740 (.CLK(clknet_leaf_19_clk),
    .D(net414),
    .RESET_B(net401),
    .Q(net500),
    .Q_N(net499));
 sky130_fd_sc_hd__dfrbp_1 merge741 (.CLK(clknet_leaf_33_clk),
    .D(net479),
    .RESET_B(net480),
    .Q(net502),
    .Q_N(net501));
 sky130_fd_sc_hd__dfrtn_1 merge742 (.CLK_N(clknet_leaf_18_clk),
    .D(net206),
    .RESET_B(net193),
    .Q(net503));
 sky130_fd_sc_hd__dfrtp_1 merge743 (.CLK(clknet_leaf_23_clk),
    .D(net448),
    .RESET_B(net451),
    .Q(net504));
 sky130_fd_sc_hd__dfrtp_1 merge744 (.CLK(clknet_leaf_21_clk),
    .D(net419),
    .RESET_B(net421),
    .Q(net505));
 sky130_fd_sc_hd__dfrtp_1 merge745 (.CLK(clknet_leaf_23_clk),
    .D(net330),
    .RESET_B(net327),
    .Q(net506));
 sky130_fd_sc_hd__dfsbp_2 merge746 (.CLK(clknet_leaf_1_clk),
    .D(net53),
    .SET_B(net55),
    .Q(net508),
    .Q_N(net507));
 sky130_fd_sc_hd__dfsbp_1 merge747 (.CLK(clknet_leaf_14_clk),
    .D(net228),
    .SET_B(net235),
    .Q(net510),
    .Q_N(net509));
 sky130_fd_sc_hd__dfstp_1 merge748 (.CLK(clknet_leaf_36_clk),
    .D(net166),
    .Q(net918));
 sky130_fd_sc_hd__dfstp_1 merge749 (.CLK(clknet_leaf_6_clk),
    .D(net139),
    .Q(net140));
 sky130_fd_sc_hd__dfstp_1 merge750 (.CLK(clknet_leaf_32_clk),
    .D(net374),
    .SET_B(net376),
    .Q(net879));
 sky130_fd_sc_hd__dlrbn_1 merge751 (.GATE_N(clknet_leaf_8_clk),
    .RESET_B(net38),
    .Q(net513),
    .Q_N(net512));
 sky130_fd_sc_hd__dlrbn_1 merge752 (.D(net82),
    .GATE_N(clknet_leaf_40_clk),
    .RESET_B(net87),
    .Q(net515),
    .Q_N(net514));
 sky130_fd_sc_hd__dlrbp_1 merge753 (.D(net60),
    .GATE(clknet_leaf_0_clk),
    .RESET_B(net66),
    .Q(net517),
    .Q_N(net516));
 sky130_fd_sc_hd__dlrbp_1 merge754 (.D(net129),
    .GATE(clknet_leaf_13_clk),
    .RESET_B(net120),
    .Q(net519),
    .Q_N(net518));
 sky130_fd_sc_hd__dlrtn_1 merge755 (.D(net259),
    .GATE_N(clknet_leaf_35_clk),
    .RESET_B(net266),
    .Q(net520));
 sky130_fd_sc_hd__dfxbp_2 s756 (.CLK(clknet_leaf_8_clk),
    .D(net30),
    .Q(net522),
    .Q_N(net521));
 sky130_fd_sc_hd__dfxbp_1 s757 (.CLK(clknet_leaf_8_clk),
    .D(net32),
    .Q(net524),
    .Q_N(net523));
 sky130_fd_sc_hd__dfxtp_4 s758 (.CLK(clknet_leaf_8_clk),
    .D(net34),
    .Q(net525));
 sky130_fd_sc_hd__dfxtp_2 s759 (.CLK(clknet_leaf_8_clk),
    .D(net35),
    .Q(net526));
 sky130_fd_sc_hd__dfxtp_2 s760 (.CLK(clknet_leaf_6_clk),
    .D(net44),
    .Q(net527));
 sky130_fd_sc_hd__dlclkp_1 s761 (.CLK(clknet_2_1__leaf_clk),
    .GATE(net45),
    .GCLK(net528));
 sky130_fd_sc_hd__dlclkp_2 s762 (.CLK(clknet_leaf_1_clk),
    .GATE(net51),
    .GCLK(net898));
 sky130_fd_sc_hd__dlclkp_4 s763 (.CLK(clknet_leaf_1_clk),
    .GATE(net58),
    .GCLK(net529));
 sky130_fd_sc_hd__dlxbn_1 s764 (.D(net63),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net933),
    .Q_N(net530));
 sky130_fd_sc_hd__dlxbn_2 s765 (.D(net65),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net532),
    .Q_N(net531));
 sky130_fd_sc_hd__dlxbp_1 s766 (.D(net68),
    .GATE(clknet_leaf_0_clk),
    .Q(net534),
    .Q_N(net533));
 sky130_fd_sc_hd__dlxtn_1 s767 (.D(net69),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net929));
 sky130_fd_sc_hd__dlxtn_2 s768 (.D(net70),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net535));
 sky130_fd_sc_hd__dlxtn_1 s769 (.D(net71),
    .GATE_N(clknet_leaf_0_clk),
    .Q(net536));
 sky130_fd_sc_hd__dlxtp_1 s770 (.D(net72),
    .GATE(clknet_leaf_0_clk),
    .Q(net537));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s771 (.D(net74),
    .SLEEP_B(clknet_leaf_0_clk),
    .Q(net930));
 sky130_fd_sc_hd__dfxbp_1 s772 (.CLK(clknet_leaf_41_clk),
    .D(net76),
    .Q(net539),
    .Q_N(net538));
 sky130_fd_sc_hd__dfxbp_1 s773 (.CLK(clknet_leaf_41_clk),
    .D(net79),
    .Q(net541),
    .Q_N(net540));
 sky130_fd_sc_hd__dfxtp_1 s774 (.CLK(clknet_leaf_41_clk),
    .D(net80),
    .Q(net914));
 sky130_fd_sc_hd__dfxtp_2 s775 (.CLK(clknet_leaf_40_clk),
    .D(net81),
    .Q(net872));
 sky130_fd_sc_hd__dfxtp_1 s776 (.CLK(clknet_leaf_40_clk),
    .D(net85),
    .Q(net887));
 sky130_fd_sc_hd__dlclkp_1 s777 (.CLK(clknet_leaf_40_clk),
    .GATE(net89),
    .GCLK(net542));
 sky130_fd_sc_hd__dlclkp_2 s778 (.CLK(clknet_leaf_9_clk),
    .GATE(net104),
    .GCLK(net543));
 sky130_fd_sc_hd__dlclkp_4 s779 (.CLK(clknet_leaf_10_clk),
    .GATE(net105),
    .GCLK(net544));
 sky130_fd_sc_hd__dlxbn_2 s780 (.D(net106),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net546),
    .Q_N(net545));
 sky130_fd_sc_hd__dlxbn_2 s781 (.D(net107),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net886),
    .Q_N(net547));
 sky130_fd_sc_hd__dlxbp_1 s782 (.D(net108),
    .GATE(clknet_leaf_10_clk),
    .Q(net549),
    .Q_N(net548));
 sky130_fd_sc_hd__dlxtn_2 s783 (.D(net109),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net550));
 sky130_fd_sc_hd__dlxtn_2 s784 (.D(net117),
    .GATE_N(clknet_leaf_9_clk),
    .Q(net551));
 sky130_fd_sc_hd__dlxtn_4 s785 (.D(net118),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net552));
 sky130_fd_sc_hd__dlxtp_1 s786 (.D(net119),
    .GATE(clknet_leaf_5_clk),
    .Q(net553));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s787 (.D(net121),
    .SLEEP_B(clknet_leaf_9_clk),
    .Q(net554));
 sky130_fd_sc_hd__dfxbp_1 s788 (.CLK(clknet_leaf_13_clk),
    .D(net123),
    .Q(net556),
    .Q_N(net555));
 sky130_fd_sc_hd__dfxbp_1 s789 (.CLK(clknet_leaf_3_clk),
    .D(net124),
    .Q(net558),
    .Q_N(net557));
 sky130_fd_sc_hd__dfxtp_2 s790 (.CLK(clknet_leaf_5_clk),
    .D(net125),
    .Q(net559));
 sky130_fd_sc_hd__dfxtp_1 s791 (.CLK(clknet_leaf_5_clk),
    .D(net126),
    .Q(net560));
 sky130_fd_sc_hd__dfxtp_4 s792 (.CLK(clknet_leaf_13_clk),
    .D(net127),
    .Q(net561));
 sky130_fd_sc_hd__dlclkp_1 s793 (.CLK(clknet_leaf_13_clk),
    .GATE(net128),
    .GCLK(net562));
 sky130_fd_sc_hd__dlclkp_2 s794 (.CLK(clknet_leaf_5_clk),
    .GATE(net130),
    .GCLK(net908));
 sky130_fd_sc_hd__dlclkp_4 s795 (.CLK(clknet_leaf_5_clk),
    .GATE(net134),
    .GCLK(net563));
 sky130_fd_sc_hd__dlxbn_2 s796 (.D(net135),
    .GATE_N(clknet_leaf_6_clk),
    .Q(net565),
    .Q_N(net564));
 sky130_fd_sc_hd__dlxbn_1 s797 (.D(net138),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net567),
    .Q_N(net566));
 sky130_fd_sc_hd__dlxbp_1 s798 (.D(net143),
    .GATE(clknet_leaf_6_clk),
    .Q(net907),
    .Q_N(net568));
 sky130_fd_sc_hd__dlxtn_4 s799 (.D(net144),
    .GATE_N(clknet_leaf_5_clk),
    .Q(net569));
 sky130_fd_sc_hd__dlxtn_2 s800 (.D(net145),
    .GATE_N(clknet_leaf_3_clk),
    .Q(net570));
 sky130_fd_sc_hd__dlxtn_2 s801 (.D(net146),
    .GATE_N(clknet_leaf_2_clk),
    .Q(net571));
 sky130_fd_sc_hd__dlxtp_1 s802 (.D(net149),
    .GATE(clknet_leaf_34_clk),
    .Q(net572));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s803 (.D(net150),
    .SLEEP_B(clknet_leaf_2_clk),
    .Q(net573));
 sky130_fd_sc_hd__dfxbp_1 s804 (.CLK(clknet_leaf_42_clk),
    .D(net151),
    .Q(net575),
    .Q_N(net574));
 sky130_fd_sc_hd__dfxbp_1 s805 (.CLK(clknet_leaf_2_clk),
    .D(net152),
    .Q(net577),
    .Q_N(net576));
 sky130_fd_sc_hd__dfxtp_4 s806 (.CLK(clknet_leaf_36_clk),
    .D(net154),
    .Q(net578));
 sky130_fd_sc_hd__dfxtp_2 s807 (.CLK(clknet_leaf_2_clk),
    .D(net155),
    .Q(net579));
 sky130_fd_sc_hd__dfxtp_1 s808 (.CLK(clknet_leaf_42_clk),
    .D(net157),
    .Q(net911));
 sky130_fd_sc_hd__dlclkp_1 s809 (.CLK(clknet_leaf_2_clk),
    .GATE(net163),
    .GCLK(net580));
 sky130_fd_sc_hd__dlclkp_2 s810 (.CLK(clknet_leaf_2_clk),
    .GATE(net168),
    .GCLK(net902));
 sky130_fd_sc_hd__dlclkp_4 s811 (.CLK(clknet_leaf_2_clk),
    .GATE(net169),
    .GCLK(net581));
 sky130_fd_sc_hd__dlxbn_1 s812 (.D(net170),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net583),
    .Q_N(net582));
 sky130_fd_sc_hd__dlxbn_1 s813 (.D(net171),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net909),
    .Q_N(net584));
 sky130_fd_sc_hd__dlxbp_1 s814 (.D(net172),
    .GATE(clknet_leaf_40_clk),
    .Q(net585));
 sky130_fd_sc_hd__dlxtn_2 s815 (.D(net173),
    .GATE_N(clknet_leaf_40_clk),
    .Q(net586));
 sky130_fd_sc_hd__dlxtn_1 s816 (.D(net174),
    .GATE_N(clknet_leaf_38_clk),
    .Q(net905));
 sky130_fd_sc_hd__dlxtn_1 s817 (.D(net175),
    .GATE_N(clknet_leaf_39_clk),
    .Q(net587));
 sky130_fd_sc_hd__dlxtp_1 s818 (.D(net179),
    .GATE(clknet_leaf_32_clk),
    .Q(net588));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s819 (.D(net180),
    .SLEEP_B(clknet_leaf_39_clk),
    .Q(net589));
 sky130_fd_sc_hd__dfxbp_1 s820 (.CLK(clknet_leaf_38_clk),
    .D(net181),
    .Q(net591),
    .Q_N(net590));
 sky130_fd_sc_hd__dfxbp_1 s821 (.CLK(clknet_leaf_38_clk),
    .D(net182),
    .Q(net593),
    .Q_N(net592));
 sky130_fd_sc_hd__dfxtp_1 s822 (.CLK(clknet_leaf_38_clk),
    .D(net183),
    .Q(net594));
 sky130_fd_sc_hd__dfxtp_1 s823 (.CLK(clknet_leaf_38_clk),
    .D(net185),
    .Q(net874));
 sky130_fd_sc_hd__dfxtp_1 s824 (.CLK(clknet_leaf_30_clk),
    .D(net186),
    .Q(net595));
 sky130_fd_sc_hd__dlclkp_1 s825 (.CLK(clknet_leaf_10_clk),
    .GATE(net198),
    .GCLK(net596));
 sky130_fd_sc_hd__dlclkp_2 s826 (.CLK(clknet_2_3__leaf_clk),
    .GATE(net199),
    .GCLK(net597));
 sky130_fd_sc_hd__dlclkp_4 s827 (.CLK(clknet_leaf_10_clk),
    .GATE(net200),
    .GCLK(net598));
 sky130_fd_sc_hd__dlxbn_2 s828 (.D(net201),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net600),
    .Q_N(net599));
 sky130_fd_sc_hd__dlxbn_1 s829 (.D(net202),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net602),
    .Q_N(net601));
 sky130_fd_sc_hd__dlxbp_1 s830 (.D(net203),
    .GATE(clknet_leaf_12_clk),
    .Q(net604),
    .Q_N(net603));
 sky130_fd_sc_hd__dlxtn_4 s831 (.D(net205),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net605));
 sky130_fd_sc_hd__dlxtn_4 s832 (.D(net209),
    .GATE_N(clknet_leaf_12_clk),
    .Q(net606));
 sky130_fd_sc_hd__dlxtn_2 s833 (.D(net210),
    .GATE_N(clknet_leaf_13_clk),
    .Q(net607));
 sky130_fd_sc_hd__dlxtp_1 s834 (.D(net212),
    .GATE(clknet_leaf_14_clk),
    .Q(net608));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s835 (.D(net213),
    .SLEEP_B(clknet_leaf_13_clk),
    .Q(net609));
 sky130_fd_sc_hd__dfxbp_2 s836 (.CLK(clknet_leaf_14_clk),
    .D(net214),
    .Q(net878),
    .Q_N(net610));
 sky130_fd_sc_hd__dfxbp_1 s837 (.CLK(clknet_leaf_14_clk),
    .D(net216),
    .Q(net612),
    .Q_N(net611));
 sky130_fd_sc_hd__dfxtp_1 s838 (.CLK(clknet_leaf_12_clk),
    .D(net217),
    .Q(net613));
 sky130_fd_sc_hd__dfxtp_4 s839 (.CLK(clknet_leaf_12_clk),
    .D(net219),
    .Q(net614));
 sky130_fd_sc_hd__dfxtp_1 s840 (.CLK(clknet_leaf_12_clk),
    .D(net221),
    .Q(net615));
 sky130_fd_sc_hd__dlclkp_1 s841 (.CLK(clknet_leaf_14_clk),
    .GATE(net223),
    .GCLK(net616));
 sky130_fd_sc_hd__dlclkp_2 s842 (.CLK(clknet_leaf_17_clk),
    .GATE(net224),
    .GCLK(net617));
 sky130_fd_sc_hd__dlclkp_4 s843 (.CLK(clknet_leaf_14_clk),
    .GATE(net225),
    .GCLK(net618));
 sky130_fd_sc_hd__dlxbn_1 s844 (.D(net227),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net620),
    .Q_N(net619));
 sky130_fd_sc_hd__dlxbn_1 s845 (.D(net231),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net622),
    .Q_N(net621));
 sky130_fd_sc_hd__dlxbp_1 s846 (.D(net232),
    .GATE(clknet_leaf_3_clk),
    .Q(net624),
    .Q_N(net623));
 sky130_fd_sc_hd__dlxtn_2 s847 (.D(net236),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net625));
 sky130_fd_sc_hd__dlxtn_1 s848 (.D(net237),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net626));
 sky130_fd_sc_hd__dlxtn_1 s849 (.D(net238),
    .GATE_N(clknet_leaf_4_clk),
    .Q(net627));
 sky130_fd_sc_hd__dlxtp_1 s850 (.D(net242),
    .GATE(clknet_leaf_4_clk),
    .Q(net628));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s851 (.D(net244),
    .SLEEP_B(clknet_leaf_15_clk),
    .Q(net629));
 sky130_fd_sc_hd__dfxbp_1 s852 (.CLK(clknet_leaf_4_clk),
    .D(net245),
    .Q(net631),
    .Q_N(net630));
 sky130_fd_sc_hd__dfxbp_2 s853 (.CLK(clknet_leaf_34_clk),
    .D(net246),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__dfxtp_1 s854 (.CLK(clknet_leaf_34_clk),
    .D(net249),
    .Q(net634));
 sky130_fd_sc_hd__dfxtp_1 s855 (.CLK(clknet_leaf_36_clk),
    .D(net250),
    .Q(net635));
 sky130_fd_sc_hd__dfxtp_1 s856 (.CLK(clknet_leaf_34_clk),
    .D(net251),
    .Q(net636));
 sky130_fd_sc_hd__dlclkp_1 s857 (.CLK(clknet_leaf_38_clk),
    .GATE(net252),
    .GCLK(net890));
 sky130_fd_sc_hd__dlclkp_2 s858 (.CLK(clknet_leaf_2_clk),
    .GATE(net256),
    .GCLK(net637));
 sky130_fd_sc_hd__dlclkp_4 s859 (.CLK(clknet_leaf_35_clk),
    .GATE(net262),
    .GCLK(net638));
 sky130_fd_sc_hd__dlxbn_2 s860 (.D(net263),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net640),
    .Q_N(net639));
 sky130_fd_sc_hd__dlxbn_1 s861 (.D(net264),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__dlxbp_1 s862 (.D(net265),
    .GATE(clknet_leaf_27_clk),
    .Q(net644),
    .Q_N(net643));
 sky130_fd_sc_hd__dlxtn_4 s863 (.D(net267),
    .GATE_N(clknet_leaf_36_clk),
    .Q(net645));
 sky130_fd_sc_hd__dlxtn_1 s864 (.D(net268),
    .GATE_N(clknet_leaf_35_clk),
    .Q(net646));
 sky130_fd_sc_hd__dlxtn_1 s865 (.D(net269),
    .GATE_N(clknet_leaf_37_clk),
    .Q(net647));
 sky130_fd_sc_hd__dlxtp_1 s866 (.D(net271),
    .GATE(clknet_leaf_38_clk),
    .Q(net648));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s867 (.D(net274),
    .SLEEP_B(clknet_leaf_36_clk),
    .Q(net649));
 sky130_fd_sc_hd__dfxbp_1 s868 (.CLK(clknet_leaf_37_clk),
    .D(net275),
    .Q(net651),
    .Q_N(net650));
 sky130_fd_sc_hd__dfxbp_1 s869 (.CLK(clknet_leaf_38_clk),
    .D(net277),
    .Q(net653),
    .Q_N(net652));
 sky130_fd_sc_hd__dfxtp_1 s870 (.CLK(clknet_leaf_37_clk),
    .D(net279),
    .Q(net654));
 sky130_fd_sc_hd__dfxtp_1 s871 (.CLK(clknet_leaf_37_clk),
    .D(net281),
    .Q(net892));
 sky130_fd_sc_hd__dfxtp_1 s872 (.CLK(clknet_leaf_37_clk),
    .D(net284),
    .Q(net655));
 sky130_fd_sc_hd__dlclkp_1 s873 (.CLK(clknet_leaf_37_clk),
    .GATE(net285),
    .GCLK(net891));
 sky130_fd_sc_hd__dlclkp_2 s874 (.CLK(clknet_leaf_37_clk),
    .GATE(net286),
    .GCLK(net656));
 sky130_fd_sc_hd__dlclkp_4 s875 (.CLK(clknet_leaf_37_clk),
    .GATE(net287),
    .GCLK(net657));
 sky130_fd_sc_hd__dlxbn_1 s876 (.D(net288),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net659),
    .Q_N(net658));
 sky130_fd_sc_hd__dlxbn_1 s877 (.D(net302),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net661),
    .Q_N(net660));
 sky130_fd_sc_hd__dlxbp_1 s878 (.D(net303),
    .GATE(clknet_leaf_19_clk),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__dlxtn_2 s879 (.D(net304),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net664));
 sky130_fd_sc_hd__dlxtn_2 s880 (.D(net305),
    .GATE_N(clknet_leaf_18_clk),
    .Q(net665));
 sky130_fd_sc_hd__dlxtn_2 s881 (.D(net306),
    .GATE_N(clknet_leaf_17_clk),
    .Q(net869));
 sky130_fd_sc_hd__dlxtp_1 s882 (.D(net311),
    .GATE(clknet_leaf_16_clk),
    .Q(net666));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s883 (.D(net315),
    .SLEEP_B(clknet_leaf_16_clk),
    .Q(net667));
 sky130_fd_sc_hd__dfxbp_1 s884 (.CLK(clknet_leaf_16_clk),
    .D(net316),
    .Q(net669),
    .Q_N(net668));
 sky130_fd_sc_hd__dfxbp_1 s885 (.CLK(clknet_leaf_23_clk),
    .D(net317),
    .Q(net671),
    .Q_N(net670));
 sky130_fd_sc_hd__dfxtp_1 s886 (.CLK(clknet_leaf_17_clk),
    .D(net318),
    .Q(net672));
 sky130_fd_sc_hd__dfxtp_2 s887 (.CLK(clknet_leaf_16_clk),
    .D(net319),
    .Q(net673));
 sky130_fd_sc_hd__dfxtp_1 s888 (.CLK(clknet_leaf_16_clk),
    .D(net320),
    .Q(net674));
 sky130_fd_sc_hd__dlclkp_1 s889 (.CLK(clknet_leaf_16_clk),
    .GATE(net323),
    .GCLK(net675));
 sky130_fd_sc_hd__dlclkp_2 s890 (.CLK(clknet_leaf_16_clk),
    .GATE(net325),
    .GCLK(net888));
 sky130_fd_sc_hd__dlclkp_4 s891 (.CLK(clknet_leaf_17_clk),
    .GATE(net326),
    .GCLK(net676));
 sky130_fd_sc_hd__dlxbn_1 s892 (.D(net328),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net678),
    .Q_N(net677));
 sky130_fd_sc_hd__dlxbn_1 s893 (.D(net334),
    .GATE_N(clknet_leaf_34_clk),
    .Q(net680),
    .Q_N(net679));
 sky130_fd_sc_hd__dlxbp_1 s894 (.D(net336),
    .GATE(clknet_leaf_15_clk),
    .Q(net682),
    .Q_N(net681));
 sky130_fd_sc_hd__dlxtn_1 s895 (.D(net338),
    .GATE_N(clknet_leaf_15_clk),
    .Q(net683));
 sky130_fd_sc_hd__dlxtn_1 s896 (.D(net341),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net684));
 sky130_fd_sc_hd__dlxtn_1 s897 (.D(net343),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net685));
 sky130_fd_sc_hd__dlxtp_1 s898 (.D(net344),
    .GATE(clknet_leaf_24_clk),
    .Q(net686));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s899 (.D(net347),
    .SLEEP_B(clknet_leaf_24_clk),
    .Q(net687));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_leaf_25_clk),
    .D(net351),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__dfxbp_1 s901 (.CLK(clknet_leaf_24_clk),
    .D(net352),
    .Q(net691),
    .Q_N(net690));
 sky130_fd_sc_hd__dfxtp_2 s902 (.CLK(clknet_leaf_24_clk),
    .D(net353),
    .Q(net692));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_leaf_31_clk),
    .D(net354),
    .Q(net693));
 sky130_fd_sc_hd__dfxtp_1 s904 (.CLK(clknet_leaf_35_clk),
    .D(net356),
    .Q(net694));
 sky130_fd_sc_hd__dlclkp_1 s905 (.CLK(clknet_leaf_26_clk),
    .GATE(net358),
    .GCLK(net695));
 sky130_fd_sc_hd__dlclkp_2 s906 (.CLK(clknet_leaf_26_clk),
    .GATE(net359),
    .GCLK(net696));
 sky130_fd_sc_hd__dlclkp_4 s907 (.CLK(clknet_leaf_34_clk),
    .GATE(net360),
    .GCLK(net697));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net361),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net698));
 sky130_fd_sc_hd__dlxbn_1 s909 (.D(net362),
    .GATE_N(clknet_leaf_32_clk),
    .Q(net699));
 sky130_fd_sc_hd__dlxbp_1 s910 (.D(net364),
    .GATE(clknet_leaf_33_clk),
    .Q(net701),
    .Q_N(net700));
 sky130_fd_sc_hd__dlxtn_1 s911 (.D(net365),
    .GATE_N(clknet_leaf_34_clk),
    .Q(net702));
 sky130_fd_sc_hd__dlxtn_1 s912 (.D(net370),
    .GATE_N(clknet_leaf_34_clk),
    .Q(net703));
 sky130_fd_sc_hd__dlxtn_1 s913 (.D(net373),
    .GATE_N(clknet_leaf_26_clk),
    .Q(net704));
 sky130_fd_sc_hd__dlxtp_1 s914 (.D(net375),
    .GATE(clknet_leaf_31_clk),
    .Q(net705));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s915 (.D(net379),
    .SLEEP_B(clknet_leaf_33_clk),
    .Q(net706));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_leaf_30_clk),
    .D(net381),
    .Q(net707));
 sky130_fd_sc_hd__dfxbp_1 s917 (.CLK(clknet_leaf_31_clk),
    .D(net383),
    .Q(net708));
 sky130_fd_sc_hd__dfxtp_1 s918 (.CLK(clknet_leaf_30_clk),
    .D(net384),
    .Q(net709));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_leaf_33_clk),
    .D(net387),
    .Q(net710));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_leaf_33_clk),
    .D(net389),
    .Q(net711));
 sky130_fd_sc_hd__dlclkp_1 s921 (.CLK(clknet_leaf_29_clk),
    .GATE(net390),
    .GCLK(net880));
 sky130_fd_sc_hd__dlclkp_2 s922 (.CLK(clknet_leaf_32_clk),
    .GATE(net393),
    .GCLK(net712));
 sky130_fd_sc_hd__dlclkp_4 s923 (.CLK(clknet_leaf_31_clk),
    .GATE(net394),
    .GCLK(net713));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net400),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net715),
    .Q_N(net714));
 sky130_fd_sc_hd__dlxbn_1 s925 (.D(net403),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net717),
    .Q_N(net716));
 sky130_fd_sc_hd__dlxbp_1 s926 (.D(net404),
    .GATE(clknet_leaf_19_clk),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dlxtn_1 s927 (.D(net406),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net720));
 sky130_fd_sc_hd__dlxtn_4 s928 (.D(net407),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net721));
 sky130_fd_sc_hd__dlxtn_2 s929 (.D(net410),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net722));
 sky130_fd_sc_hd__dlxtp_1 s930 (.D(net412),
    .GATE(clknet_leaf_19_clk),
    .Q(net723));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s931 (.D(net413),
    .SLEEP_B(clknet_leaf_20_clk),
    .Q(net724));
 sky130_fd_sc_hd__dfxbp_1 s932 (.CLK(clknet_leaf_21_clk),
    .D(net420),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__dfxbp_1 s933 (.CLK(clknet_leaf_21_clk),
    .D(net423),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dfxtp_2 s934 (.CLK(clknet_leaf_21_clk),
    .D(net424),
    .Q(net729));
 sky130_fd_sc_hd__dfxtp_2 s935 (.CLK(clknet_leaf_21_clk),
    .D(net425),
    .Q(net730));
 sky130_fd_sc_hd__dfxtp_2 s936 (.CLK(clknet_leaf_21_clk),
    .D(net426),
    .Q(net731));
 sky130_fd_sc_hd__dlclkp_1 s937 (.CLK(clknet_leaf_22_clk),
    .GATE(net430),
    .GCLK(net732));
 sky130_fd_sc_hd__dlclkp_2 s938 (.CLK(clknet_leaf_23_clk),
    .GATE(net431),
    .GCLK(net733));
 sky130_fd_sc_hd__dlclkp_4 s939 (.CLK(clknet_leaf_22_clk),
    .GATE(net432),
    .GCLK(net734));
 sky130_fd_sc_hd__dlxbn_1 s940 (.D(net433),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__dlxbn_1 s941 (.D(net434),
    .GATE_N(clknet_leaf_23_clk),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__dlxbp_1 s942 (.D(net435),
    .GATE(clknet_leaf_21_clk),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__dlxtn_1 s943 (.D(net436),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net741));
 sky130_fd_sc_hd__dlxtn_1 s944 (.D(net437),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net742));
 sky130_fd_sc_hd__dlxtn_1 s945 (.D(net438),
    .GATE_N(clknet_leaf_22_clk),
    .Q(net743));
 sky130_fd_sc_hd__dlxtp_1 s946 (.D(net445),
    .GATE(clknet_leaf_24_clk),
    .Q(net744));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s947 (.D(net447),
    .SLEEP_B(clknet_leaf_22_clk),
    .Q(net745));
 sky130_fd_sc_hd__dfxbp_1 s948 (.CLK(clknet_leaf_28_clk),
    .D(net455),
    .Q(net746));
 sky130_fd_sc_hd__dfxbp_1 s949 (.CLK(clknet_leaf_27_clk),
    .D(net456),
    .Q(net748),
    .Q_N(net747));
 sky130_fd_sc_hd__dfxtp_1 s950 (.CLK(clknet_leaf_29_clk),
    .D(net458),
    .Q(net749));
 sky130_fd_sc_hd__dfxtp_1 s951 (.CLK(clknet_leaf_28_clk),
    .D(net459),
    .Q(net750));
 sky130_fd_sc_hd__dfxtp_1 s952 (.CLK(clknet_leaf_27_clk),
    .D(net460),
    .Q(net751));
 sky130_fd_sc_hd__dlclkp_1 s953 (.CLK(clknet_leaf_26_clk),
    .GATE(net461),
    .GCLK(net752));
 sky130_fd_sc_hd__dlclkp_2 s954 (.CLK(clknet_leaf_28_clk),
    .GATE(net462),
    .GCLK(net753));
 sky130_fd_sc_hd__dlclkp_4 s955 (.CLK(clknet_leaf_28_clk),
    .GATE(net466),
    .GCLK(net754));
 sky130_fd_sc_hd__dlxbn_1 s956 (.D(net468),
    .GATE_N(clknet_leaf_28_clk),
    .Q(net755));
 sky130_fd_sc_hd__dlxbn_1 s957 (.D(net469),
    .GATE_N(clknet_leaf_30_clk),
    .Q(net756));
 sky130_fd_sc_hd__dlxbp_1 s958 (.D(net470),
    .GATE(clknet_leaf_30_clk),
    .Q(net758),
    .Q_N(net757));
 sky130_fd_sc_hd__dlxtn_1 s959 (.D(net475),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net759));
 sky130_fd_sc_hd__dlxtn_1 s960 (.D(net477),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net760));
 sky130_fd_sc_hd__dlxtn_1 s961 (.D(net478),
    .GATE_N(clknet_leaf_29_clk),
    .Q(net761));
 sky130_fd_sc_hd__dlxtp_1 s962 (.D(net481),
    .GATE(clknet_leaf_30_clk),
    .Q(net762));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s963 (.D(net483),
    .SLEEP_B(clknet_leaf_27_clk),
    .Q(net763));
 sky130_fd_sc_hd__dfxbp_1 s964 (.CLK(clknet_leaf_30_clk),
    .D(net485),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dfxbp_1 s965 (.CLK(clknet_leaf_30_clk),
    .D(net486),
    .Q(net766));
 sky130_fd_sc_hd__dfxtp_1 s966 (.CLK(clknet_leaf_30_clk),
    .D(net489),
    .Q(net767));
 sky130_fd_sc_hd__dfxtp_1 s967 (.CLK(clknet_leaf_29_clk),
    .D(net491),
    .Q(net768));
 sky130_fd_sc_hd__dfxtp_1 s968 (.CLK(clknet_leaf_33_clk),
    .D(net494),
    .Q(net769));
 sky130_fd_sc_hd__dlclkp_1 s969 (.CLK(clknet_leaf_30_clk),
    .GATE(net497),
    .GCLK(net770));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in0),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(in1),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net771));
 sky130_fd_sc_hd__buf_2 input4 (.A(in11),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in12),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(in13),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in14),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input8 (.A(in15),
    .X(net776));
 sky130_fd_sc_hd__buf_2 input9 (.A(in16),
    .X(net777));
 sky130_fd_sc_hd__buf_2 input10 (.A(in17),
    .X(net778));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(in18),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in19),
    .X(net780));
 sky130_fd_sc_hd__buf_2 input13 (.A(in2),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in20),
    .X(net782));
 sky130_fd_sc_hd__buf_2 input15 (.A(in21),
    .X(net783));
 sky130_fd_sc_hd__buf_2 input16 (.A(in22),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in23),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in25),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(in26),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in27),
    .X(net789));
 sky130_fd_sc_hd__buf_4 input22 (.A(in28),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_8 input23 (.A(in29),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(in3),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in30),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in31),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in32),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(in33),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(in34),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in35),
    .X(net798));
 sky130_fd_sc_hd__buf_4 input31 (.A(in36),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(in37),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(in38),
    .X(net801));
 sky130_fd_sc_hd__buf_4 input34 (.A(in39),
    .X(net802));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(in4),
    .X(net803));
 sky130_fd_sc_hd__buf_2 input36 (.A(in40),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in41),
    .X(net805));
 sky130_fd_sc_hd__buf_1 input38 (.A(in42),
    .X(net806));
 sky130_fd_sc_hd__buf_2 input39 (.A(in43),
    .X(net807));
 sky130_fd_sc_hd__buf_2 input40 (.A(in44),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in45),
    .X(net809));
 sky130_fd_sc_hd__buf_1 input42 (.A(in46),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in47),
    .X(net811));
 sky130_fd_sc_hd__buf_1 input44 (.A(in48),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(in49),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in5),
    .X(net814));
 sky130_fd_sc_hd__buf_2 input47 (.A(in50),
    .X(net815));
 sky130_fd_sc_hd__buf_4 input48 (.A(in51),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(in52),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(in53),
    .X(net818));
 sky130_fd_sc_hd__buf_4 input51 (.A(in54),
    .X(net819));
 sky130_fd_sc_hd__buf_1 input52 (.A(in55),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in56),
    .X(net821));
 sky130_fd_sc_hd__buf_1 input54 (.A(in57),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in58),
    .X(net823));
 sky130_fd_sc_hd__buf_1 input56 (.A(in59),
    .X(net824));
 sky130_fd_sc_hd__buf_1 input57 (.A(in6),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(in60),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(in61),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in62),
    .X(net828));
 sky130_fd_sc_hd__buf_1 input61 (.A(in63),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(in64),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(in65),
    .X(net831));
 sky130_fd_sc_hd__buf_1 input64 (.A(in66),
    .X(net832));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(in67),
    .X(net833));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(in68),
    .X(net834));
 sky130_fd_sc_hd__buf_2 input67 (.A(in69),
    .X(net835));
 sky130_fd_sc_hd__buf_6 input68 (.A(in7),
    .X(net836));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(in70),
    .X(net837));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(in71),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(in72),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(in73),
    .X(net840));
 sky130_fd_sc_hd__buf_2 input73 (.A(in74),
    .X(net841));
 sky130_fd_sc_hd__buf_1 input74 (.A(in75),
    .X(net842));
 sky130_fd_sc_hd__buf_1 input75 (.A(in76),
    .X(net843));
 sky130_fd_sc_hd__buf_4 input76 (.A(in77),
    .X(net844));
 sky130_fd_sc_hd__buf_1 input77 (.A(in78),
    .X(net845));
 sky130_fd_sc_hd__buf_1 input78 (.A(in79),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(in8),
    .X(net847));
 sky130_fd_sc_hd__buf_1 input80 (.A(in80),
    .X(net848));
 sky130_fd_sc_hd__buf_1 input81 (.A(in81),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(in82),
    .X(net850));
 sky130_fd_sc_hd__buf_1 input83 (.A(in83),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(in84),
    .X(net852));
 sky130_fd_sc_hd__buf_1 input85 (.A(in85),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(in86),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(in87),
    .X(net855));
 sky130_fd_sc_hd__buf_1 input88 (.A(in88),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(in89),
    .X(net857));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(in9),
    .X(net858));
 sky130_fd_sc_hd__buf_1 input91 (.A(in90),
    .X(net859));
 sky130_fd_sc_hd__buf_2 input92 (.A(in91),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(in92),
    .X(net861));
 sky130_fd_sc_hd__buf_1 input94 (.A(in93),
    .X(net862));
 sky130_fd_sc_hd__buf_1 input95 (.A(in94),
    .X(net863));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(in95),
    .X(net864));
 sky130_fd_sc_hd__buf_1 input97 (.A(in96),
    .X(net865));
 sky130_fd_sc_hd__buf_2 input98 (.A(in97),
    .X(net866));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(in98),
    .X(net867));
 sky130_fd_sc_hd__dlymetal6s2s_1 input100 (.A(in99),
    .X(net868));
 sky130_fd_sc_hd__buf_2 output101 (.A(net869),
    .X(out0));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(clknet_1_0__leaf_net870),
    .X(out1));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net871),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output104 (.A(net872),
    .X(out11));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net873),
    .X(out12));
 sky130_fd_sc_hd__buf_2 output106 (.A(net874),
    .X(out13));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net957),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output108 (.A(net876),
    .X(out15));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net877),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output110 (.A(net878),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output111 (.A(net879),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net880),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net881),
    .X(out21));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(clknet_1_1__leaf_net882),
    .X(out22));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(clknet_1_0__leaf_net883),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(clknet_1_0__leaf_net884),
    .X(out26));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(clknet_1_0__leaf_net885),
    .X(out27));
 sky130_fd_sc_hd__buf_2 output118 (.A(net886),
    .X(out28));
 sky130_fd_sc_hd__buf_2 output119 (.A(net887),
    .X(out29));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(clknet_1_0__leaf_net888),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output121 (.A(net889),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(clknet_1_1__leaf_net890),
    .X(out31));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net891),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output124 (.A(net892),
    .X(out34));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(clknet_1_0__leaf_net893),
    .X(out35));
 sky130_fd_sc_hd__buf_2 output126 (.A(net944),
    .X(out37));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net895),
    .X(out38));
 sky130_fd_sc_hd__buf_2 output128 (.A(net896),
    .X(out4));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(clknet_1_1__leaf_net897),
    .X(out41));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(clknet_1_0__leaf_net898),
    .X(out42));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(clknet_1_0__leaf_net899),
    .X(out43));
 sky130_fd_sc_hd__buf_2 output132 (.A(net900),
    .X(out44));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net901),
    .X(out45));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(clknet_1_0__leaf_net902),
    .X(out46));
 sky130_fd_sc_hd__buf_4 output135 (.A(net903),
    .X(out47));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(clknet_1_1__leaf_net904),
    .X(out49));
 sky130_fd_sc_hd__buf_2 output137 (.A(net905),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output138 (.A(net906),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output139 (.A(net907),
    .X(out51));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(clknet_1_0__leaf_net908),
    .X(out52));
 sky130_fd_sc_hd__buf_2 output141 (.A(net909),
    .X(out54));
 sky130_fd_sc_hd__buf_2 output142 (.A(net910),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output143 (.A(net911),
    .X(out57));
 sky130_fd_sc_hd__buf_2 output144 (.A(net912),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output145 (.A(net913),
    .X(out59));
 sky130_fd_sc_hd__buf_2 output146 (.A(net914),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output147 (.A(net949),
    .X(out60));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(clknet_1_1__leaf_net916),
    .X(out61));
 sky130_fd_sc_hd__buf_2 output149 (.A(net917),
    .X(out62));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(clknet_1_0__leaf_net918),
    .X(out63));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net919),
    .X(out65));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(clknet_1_0__leaf_net920),
    .X(out67));
 sky130_fd_sc_hd__buf_2 output153 (.A(net921),
    .X(out68));
 sky130_fd_sc_hd__buf_2 output154 (.A(net922),
    .X(out69));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(clknet_1_0__leaf_net923),
    .X(out70));
 sky130_fd_sc_hd__buf_2 output156 (.A(net924),
    .X(out71));
 sky130_fd_sc_hd__buf_2 output157 (.A(net925),
    .X(out73));
 sky130_fd_sc_hd__buf_2 output158 (.A(net926),
    .X(out75));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(clknet_1_0__leaf_net927),
    .X(out78));
 sky130_fd_sc_hd__buf_2 output160 (.A(net928),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output161 (.A(net929),
    .X(out82));
 sky130_fd_sc_hd__buf_2 output162 (.A(net930),
    .X(out83));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(clknet_1_0__leaf_net931),
    .X(out84));
 sky130_fd_sc_hd__buf_2 output164 (.A(net1068),
    .X(out85));
 sky130_fd_sc_hd__buf_2 output165 (.A(net933),
    .X(out86));
 sky130_fd_sc_hd__buf_2 output166 (.A(net934),
    .X(out88));
 sky130_fd_sc_hd__buf_2 output167 (.A(net935),
    .X(out89));
 sky130_fd_sc_hd__buf_2 output168 (.A(net936),
    .X(out90));
 sky130_fd_sc_hd__buf_2 output169 (.A(net937),
    .X(out92));
 sky130_fd_sc_hd__buf_2 output170 (.A(net938),
    .X(out94));
 sky130_fd_sc_hd__buf_2 output171 (.A(net939),
    .X(out97));
 sky130_fd_sc_hd__buf_2 output172 (.A(net940),
    .X(out99));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net67),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net197),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net37),
    .X(net943));
 sky130_fd_sc_hd__buf_12 fanout176 (.A(net894),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net191),
    .X(net945));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net36),
    .X(net946));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net36),
    .X(net947));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(net29),
    .X(net948));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net915),
    .X(net949));
 sky130_fd_sc_hd__buf_8 fanout182 (.A(net24),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(net19),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(net92),
    .X(net953));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net957),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net875),
    .X(net957));
 sky130_fd_sc_hd__buf_8 fanout190 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__buf_12 fanout192 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__buf_8 fanout193 (.A(net16),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net14),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net14),
    .X(net963));
 sky130_fd_sc_hd__buf_8 fanout196 (.A(net12),
    .X(net964));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net11),
    .X(net965));
 sky130_fd_sc_hd__buf_12 fanout198 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_8 fanout200 (.A(net10),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net912),
    .X(net969));
 sky130_fd_sc_hd__buf_12 fanout202 (.A(net9),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net22),
    .X(net972));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(net8),
    .X(net973));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(net8),
    .X(net974));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net7),
    .X(net975));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(net6),
    .X(net976));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net26),
    .X(net977));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(net921),
    .X(net978));
 sky130_fd_sc_hd__buf_2 fanout211 (.A(net5),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net550),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_2 fanout213 (.A(net550),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net550),
    .X(net982));
 sky130_fd_sc_hd__buf_8 fanout215 (.A(net4),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(net858),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net777),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net848),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net989),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net776),
    .X(net989));
 sky130_fd_sc_hd__buf_8 fanout222 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__buf_12 fanout223 (.A(net847),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net847),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net775),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net775),
    .X(net995));
 sky130_fd_sc_hd__buf_12 fanout228 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_12 fanout229 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__buf_12 fanout230 (.A(net836),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net774),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net825),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net773),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net773),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net815),
    .X(net1003));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout236 (.A(net815),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(net772),
    .X(net1005));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net805),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net805),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_8 fanout240 (.A(net803),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net801),
    .X(net1009));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net798),
    .X(net1010));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net771),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net785),
    .X(net1013));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net782),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_8 fanout247 (.A(net781),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout248 (.A(net780),
    .X(net1016));
 sky130_fd_sc_hd__buf_2 fanout249 (.A(net780),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout250 (.A(net779),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net39),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net754 (.A(net754),
    .X(clknet_0_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net754 (.A(clknet_0_net754),
    .X(clknet_1_0__leaf_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net754 (.A(clknet_0_net754),
    .X(clknet_1_1__leaf_net754));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net467 (.A(net467),
    .X(clknet_0_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_0__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net467 (.A(clknet_0_net467),
    .X(clknet_1_1__leaf_net467));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net753 (.A(net753),
    .X(clknet_0_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_0__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net753 (.A(clknet_0_net753),
    .X(clknet_1_1__leaf_net753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net752 (.A(net752),
    .X(clknet_0_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_0__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net752 (.A(clknet_0_net752),
    .X(clknet_1_1__leaf_net752));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net734 (.A(net734),
    .X(clknet_0_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_0__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net734 (.A(clknet_0_net734),
    .X(clknet_1_1__leaf_net734));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net733 (.A(net733),
    .X(clknet_0_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_0__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net733 (.A(clknet_0_net733),
    .X(clknet_1_1__leaf_net733));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net732 (.A(net732),
    .X(clknet_0_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net732 (.A(clknet_0_net732),
    .X(clknet_1_0__leaf_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net732 (.A(clknet_0_net732),
    .X(clknet_1_1__leaf_net732));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net452 (.A(net452),
    .X(clknet_0_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_0__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net452 (.A(clknet_0_net452),
    .X(clknet_1_1__leaf_net452));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net476 (.A(net476),
    .X(clknet_0_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_0__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net476 (.A(clknet_0_net476),
    .X(clknet_1_1__leaf_net476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net446 (.A(net446),
    .X(clknet_0_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_0__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net446 (.A(clknet_0_net446),
    .X(clknet_1_1__leaf_net446));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net696 (.A(net696),
    .X(clknet_0_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_0__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_1__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net676 (.A(net676),
    .X(clknet_0_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_0__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net676 (.A(clknet_0_net676),
    .X(clknet_1_1__leaf_net676));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net417 (.A(net417),
    .X(clknet_0_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_0__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net417 (.A(clknet_0_net417),
    .X(clknet_1_1__leaf_net417));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net416 (.A(net416),
    .X(clknet_0_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_0__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net416 (.A(clknet_0_net416),
    .X(clknet_1_1__leaf_net416));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net346 (.A(net346),
    .X(clknet_0_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_0__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net346 (.A(clknet_0_net346),
    .X(clknet_1_1__leaf_net346));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net349 (.A(net349),
    .X(clknet_0_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_0__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net349 (.A(clknet_0_net349),
    .X(clknet_1_1__leaf_net349));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net339 (.A(net339),
    .X(clknet_0_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_0__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_1__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net348 (.A(net348),
    .X(clknet_0_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_0__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net348 (.A(clknet_0_net348),
    .X(clknet_1_1__leaf_net348));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net888 (.A(net888),
    .X(clknet_0_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net888 (.A(clknet_0_net888),
    .X(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net444 (.A(net444),
    .X(clknet_0_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_0__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net444 (.A(clknet_0_net444),
    .X(clknet_1_1__leaf_net444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net428 (.A(net428),
    .X(clknet_0_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_0__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net428 (.A(clknet_0_net428),
    .X(clknet_1_1__leaf_net428));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net418 (.A(net418),
    .X(clknet_0_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_0__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net418 (.A(clknet_0_net418),
    .X(clknet_1_1__leaf_net418));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net367 (.A(net367),
    .X(clknet_0_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_0__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net367 (.A(clknet_0_net367),
    .X(clknet_1_1__leaf_net367));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net372 (.A(net372),
    .X(clknet_0_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_0__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net372 (.A(clknet_0_net372),
    .X(clknet_1_1__leaf_net372));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net675 (.A(net675),
    .X(clknet_0_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_0__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net675 (.A(clknet_0_net675),
    .X(clknet_1_1__leaf_net675));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net324 (.A(net324),
    .X(clknet_0_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_0__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net324 (.A(clknet_0_net324),
    .X(clknet_1_1__leaf_net324));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net638 (.A(net638),
    .X(clknet_0_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_0__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net638 (.A(clknet_0_net638),
    .X(clknet_1_1__leaf_net638));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net357 (.A(net357),
    .X(clknet_0_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_0__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net357 (.A(clknet_0_net357),
    .X(clknet_1_1__leaf_net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net637 (.A(net637),
    .X(clknet_0_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_0__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net637 (.A(clknet_0_net637),
    .X(clknet_1_1__leaf_net637));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net261 (.A(net261),
    .X(clknet_0_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_0__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net261 (.A(clknet_0_net261),
    .X(clknet_1_1__leaf_net261));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net258 (.A(net258),
    .X(clknet_0_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_0__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net258 (.A(clknet_0_net258),
    .X(clknet_1_1__leaf_net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net257 (.A(net257),
    .X(clknet_0_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_0__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net257 (.A(clknet_0_net257),
    .X(clknet_1_1__leaf_net257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net890 (.A(net890),
    .X(clknet_0_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_0__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net890 (.A(clknet_0_net890),
    .X(clknet_1_1__leaf_net890));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net618 (.A(net618),
    .X(clknet_0_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_0__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net618 (.A(clknet_0_net618),
    .X(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net388 (.A(net388),
    .X(clknet_0_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_0__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net388 (.A(clknet_0_net388),
    .X(clknet_1_1__leaf_net388));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net617 (.A(net617),
    .X(clknet_0_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_0__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net617 (.A(clknet_0_net617),
    .X(clknet_1_1__leaf_net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net313 (.A(net313),
    .X(clknet_0_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_0__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net616 (.A(net616),
    .X(clknet_0_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_0__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net616 (.A(clknet_0_net616),
    .X(clknet_1_1__leaf_net616));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net598 (.A(net598),
    .X(clknet_0_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_0__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net598 (.A(clknet_0_net598),
    .X(clknet_1_1__leaf_net598));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net241 (.A(net241),
    .X(clknet_0_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_0__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net241 (.A(clknet_0_net241),
    .X(clknet_1_1__leaf_net241));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net240 (.A(net240),
    .X(clknet_0_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_0__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net240 (.A(clknet_0_net240),
    .X(clknet_1_1__leaf_net240));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net329 (.A(net329),
    .X(clknet_0_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_0__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net329 (.A(clknet_0_net329),
    .X(clknet_1_1__leaf_net329));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net204 (.A(net204),
    .X(clknet_0_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net204 (.A(clknet_0_net204),
    .X(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net411 (.A(net411),
    .X(clknet_0_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_0__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net411 (.A(clknet_0_net411),
    .X(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net399 (.A(net399),
    .X(clknet_0_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_0__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net399 (.A(clknet_0_net399),
    .X(clknet_1_1__leaf_net399));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net340 (.A(net340),
    .X(clknet_0_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_0__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net340 (.A(clknet_0_net340),
    .X(clknet_1_1__leaf_net340));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net312 (.A(net312),
    .X(clknet_0_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_0__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net312 (.A(clknet_0_net312),
    .X(clknet_1_1__leaf_net312));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net581 (.A(net581),
    .X(clknet_0_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_0__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net581 (.A(clknet_0_net581),
    .X(clknet_1_1__leaf_net581));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net580 (.A(net580),
    .X(clknet_0_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_0__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net580 (.A(clknet_0_net580),
    .X(clknet_1_1__leaf_net580));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net918 (.A(net918),
    .X(clknet_0_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_0__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net918 (.A(clknet_0_net918),
    .X(clknet_1_1__leaf_net918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net563 (.A(net563),
    .X(clknet_0_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_0__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net563 (.A(clknet_0_net563),
    .X(clknet_1_1__leaf_net563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net247 (.A(net247),
    .X(clknet_0_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_0__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net247 (.A(clknet_0_net247),
    .X(clknet_1_1__leaf_net247));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net148 (.A(net148),
    .X(clknet_0_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_0__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net148 (.A(clknet_0_net148),
    .X(clknet_1_1__leaf_net148));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net884 (.A(net884),
    .X(clknet_0_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net884 (.A(clknet_0_net884),
    .X(clknet_1_1__leaf_net884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net229 (.A(net229),
    .X(clknet_0_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_0__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net229 (.A(clknet_0_net229),
    .X(clknet_1_1__leaf_net229));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net337 (.A(net337),
    .X(clknet_0_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_0__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net337 (.A(clknet_0_net337),
    .X(clknet_1_1__leaf_net337));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net342 (.A(net342),
    .X(clknet_0_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_0__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net342 (.A(clknet_0_net342),
    .X(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net893 (.A(net893),
    .X(clknet_0_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_0__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net893 (.A(clknet_0_net893),
    .X(clknet_1_1__leaf_net893));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net280 (.A(net280),
    .X(clknet_0_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_0__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net280 (.A(clknet_0_net280),
    .X(clknet_1_1__leaf_net280));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net282 (.A(net282),
    .X(clknet_0_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_0__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net282 (.A(clknet_0_net282),
    .X(clknet_1_1__leaf_net282));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net141 (.A(net141),
    .X(clknet_0_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_0__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_1__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net147 (.A(net147),
    .X(clknet_0_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_0__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net147 (.A(clknet_0_net147),
    .X(clknet_1_1__leaf_net147));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net156 (.A(net156),
    .X(clknet_0_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_0__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net156 (.A(clknet_0_net156),
    .X(clknet_1_1__leaf_net156));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net159 (.A(net159),
    .X(clknet_0_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_0__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net159 (.A(clknet_0_net159),
    .X(clknet_1_1__leaf_net159));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net908 (.A(net908),
    .X(clknet_0_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_0__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net908 (.A(clknet_0_net908),
    .X(clknet_1_1__leaf_net908));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net870 (.A(net870),
    .X(clknet_0_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net870 (.A(clknet_0_net870),
    .X(clknet_1_0__leaf_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net870 (.A(clknet_0_net870),
    .X(clknet_1_1__leaf_net870));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net136 (.A(net136),
    .X(clknet_0_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_0__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net136 (.A(clknet_0_net136),
    .X(clknet_1_1__leaf_net136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net544 (.A(net544),
    .X(clknet_0_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net544 (.A(clknet_0_net544),
    .X(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net363 (.A(net363),
    .X(clknet_0_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_0__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net363 (.A(clknet_0_net363),
    .X(clknet_1_1__leaf_net363));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net291 (.A(net291),
    .X(clknet_0_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net291 (.A(clknet_0_net291),
    .X(clknet_1_1__leaf_net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net405 (.A(net405),
    .X(clknet_0_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_0__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net405 (.A(clknet_0_net405),
    .X(clknet_1_1__leaf_net405));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net397 (.A(net397),
    .X(clknet_0_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_0__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net397 (.A(clknet_0_net397),
    .X(clknet_1_1__leaf_net397));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net415 (.A(net415),
    .X(clknet_0_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_0__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_1__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net409 (.A(net409),
    .X(clknet_0_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_0__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net409 (.A(clknet_0_net409),
    .X(clknet_1_1__leaf_net409));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net396 (.A(net396),
    .X(clknet_0_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_0__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net396 (.A(clknet_0_net396),
    .X(clknet_1_1__leaf_net396));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net408 (.A(net408),
    .X(clknet_0_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_0__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net408 (.A(clknet_0_net408),
    .X(clknet_1_1__leaf_net408));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net297 (.A(net297),
    .X(clknet_0_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_0__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_1__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net299 (.A(net299),
    .X(clknet_0_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net299 (.A(clknet_0_net299),
    .X(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net295 (.A(net295),
    .X(clknet_0_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_0__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net295 (.A(clknet_0_net295),
    .X(clknet_1_1__leaf_net295));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net131 (.A(net131),
    .X(clknet_0_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_0__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_1__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net132 (.A(net132),
    .X(clknet_0_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_0__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net132 (.A(clknet_0_net132),
    .X(clknet_1_1__leaf_net132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net883 (.A(net883),
    .X(clknet_0_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net883 (.A(clknet_0_net883),
    .X(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net112 (.A(net112),
    .X(clknet_0_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_0__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net112 (.A(clknet_0_net112),
    .X(clknet_1_1__leaf_net112));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net114 (.A(net114),
    .X(clknet_0_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_0__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net114 (.A(clknet_0_net114),
    .X(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net133 (.A(net133),
    .X(clknet_0_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net133 (.A(clknet_0_net133),
    .X(clknet_1_1__leaf_net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net899 (.A(net899),
    .X(clknet_0_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_0__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net899 (.A(clknet_0_net899),
    .X(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net116 (.A(net116),
    .X(clknet_0_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_0__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net116 (.A(clknet_0_net116),
    .X(clknet_1_1__leaf_net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net122 (.A(net122),
    .X(clknet_0_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_0__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net122 (.A(clknet_0_net122),
    .X(clknet_1_1__leaf_net122));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net115 (.A(net115),
    .X(clknet_0_net115));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net115 (.A(clknet_0_net115),
    .X(clknet_1_0__leaf_net115));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net115 (.A(clknet_0_net115),
    .X(clknet_1_1__leaf_net115));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net278 (.A(net278),
    .X(clknet_0_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_0__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net278 (.A(clknet_0_net278),
    .X(clknet_1_1__leaf_net278));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net543 (.A(net543),
    .X(clknet_0_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net543 (.A(clknet_0_net543),
    .X(clknet_1_0__leaf_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net543 (.A(clknet_0_net543),
    .X(clknet_1_1__leaf_net543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net207 (.A(net207),
    .X(clknet_0_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_0__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net207 (.A(clknet_0_net207),
    .X(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net429 (.A(net429),
    .X(clknet_0_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_0__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net429 (.A(clknet_0_net429),
    .X(clknet_1_1__leaf_net429));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net220 (.A(net220),
    .X(clknet_0_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net220 (.A(clknet_0_net220),
    .X(clknet_1_1__leaf_net220));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net194 (.A(net194),
    .X(clknet_0_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_0__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net194 (.A(clknet_0_net194),
    .X(clknet_1_1__leaf_net194));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net111 (.A(net111),
    .X(clknet_0_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_0__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net111 (.A(clknet_0_net111),
    .X(clknet_1_1__leaf_net111));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net542 (.A(net542),
    .X(clknet_0_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_0__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net542 (.A(clknet_0_net542),
    .X(clknet_1_1__leaf_net542));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net529 (.A(net529),
    .X(clknet_0_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_0__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net529 (.A(clknet_0_net529),
    .X(clknet_1_1__leaf_net529));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net904 (.A(net904),
    .X(clknet_0_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_0__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net904 (.A(clknet_0_net904),
    .X(clknet_1_1__leaf_net904));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net885 (.A(net885),
    .X(clknet_0_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_0__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net885 (.A(clknet_0_net885),
    .X(clknet_1_1__leaf_net885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net83 (.A(net83),
    .X(clknet_0_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_0__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net83 (.A(clknet_0_net83),
    .X(clknet_1_1__leaf_net83));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net56 (.A(net56),
    .X(clknet_0_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net56 (.A(clknet_0_net56),
    .X(clknet_1_0__leaf_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net56 (.A(clknet_0_net56),
    .X(clknet_1_1__leaf_net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net62 (.A(net62),
    .X(clknet_0_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net62 (.A(clknet_0_net62),
    .X(clknet_1_0__leaf_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net62 (.A(clknet_0_net62),
    .X(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net59 (.A(net59),
    .X(clknet_0_net59));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net59 (.A(clknet_0_net59),
    .X(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net59 (.A(clknet_0_net59),
    .X(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net254 (.A(net254),
    .X(clknet_0_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_0__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net254 (.A(clknet_0_net254),
    .X(clknet_1_1__leaf_net254));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net253 (.A(net253),
    .X(clknet_0_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_0__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net253 (.A(clknet_0_net253),
    .X(clknet_1_1__leaf_net253));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net248 (.A(net248),
    .X(clknet_0_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_0__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net248 (.A(clknet_0_net248),
    .X(clknet_1_1__leaf_net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net920 (.A(net920),
    .X(clknet_0_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_0__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net920 (.A(clknet_0_net920),
    .X(clknet_1_1__leaf_net920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net927 (.A(net927),
    .X(clknet_0_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_0__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net927 (.A(clknet_0_net927),
    .X(clknet_1_1__leaf_net927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net64 (.A(net64),
    .X(clknet_0_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net64 (.A(clknet_0_net64),
    .X(clknet_1_0__leaf_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net64 (.A(clknet_0_net64),
    .X(clknet_1_1__leaf_net64));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net61 (.A(net61),
    .X(clknet_0_net61));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net61 (.A(clknet_0_net61),
    .X(clknet_1_0__leaf_net61));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net61 (.A(clknet_0_net61),
    .X(clknet_1_1__leaf_net61));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net57 (.A(net57),
    .X(clknet_0_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net57 (.A(clknet_0_net57),
    .X(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net57 (.A(clknet_0_net57),
    .X(clknet_1_1__leaf_net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net78 (.A(net78),
    .X(clknet_0_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_0__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net78 (.A(clknet_0_net78),
    .X(clknet_1_1__leaf_net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net923 (.A(net923),
    .X(clknet_0_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net75 (.A(net75),
    .X(clknet_0_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_0__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net75 (.A(clknet_0_net75),
    .X(clknet_1_1__leaf_net75));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net916 (.A(net916),
    .X(clknet_0_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_0__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net916 (.A(clknet_0_net916),
    .X(clknet_1_1__leaf_net916));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net528 (.A(net528),
    .X(clknet_0_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net158 (.A(net158),
    .X(clknet_0_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_0__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net158 (.A(clknet_0_net158),
    .X(clknet_1_1__leaf_net158));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net160 (.A(net160),
    .X(clknet_0_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_0__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net160 (.A(clknet_0_net160),
    .X(clknet_1_1__leaf_net160));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net47 (.A(net47),
    .X(clknet_0_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net47 (.A(clknet_0_net47),
    .X(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net47 (.A(clknet_0_net47),
    .X(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net882 (.A(net882),
    .X(clknet_0_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net243 (.A(net243),
    .X(clknet_0_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_0__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net243 (.A(clknet_0_net243),
    .X(clknet_1_1__leaf_net243));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net73 (.A(net73),
    .X(clknet_0_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net73 (.A(clknet_0_net73),
    .X(clknet_1_0__leaf_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net73 (.A(clknet_0_net73),
    .X(clknet_1_1__leaf_net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net54 (.A(net54),
    .X(clknet_0_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_0__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net54 (.A(clknet_0_net54),
    .X(clknet_1_1__leaf_net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net137 (.A(net137),
    .X(clknet_0_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_0__leaf_net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net137 (.A(clknet_0_net137),
    .X(clknet_1_1__leaf_net137));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(net1031),
    .X(net1020));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net987),
    .A1(net13),
    .A2(net966),
    .A3(net1016),
    .S0(net1056),
    .S1(net1101),
    .X(net1021));
 sky130_fd_sc_hd__mux4_1 clone3 (.A0(net1070),
    .A1(net794),
    .A2(net1024),
    .A3(net27),
    .S0(net1026),
    .S1(net971),
    .X(net1022));
 sky130_fd_sc_hd__mux4_1 clone4 (.A0(net969),
    .A1(net1026),
    .A2(net1059),
    .A3(net932),
    .S0(net1070),
    .S1(net985),
    .X(net1023));
 sky130_fd_sc_hd__mux4_1 clone5 (.A0(net976),
    .A1(net964),
    .A2(net1056),
    .A3(net965),
    .S0(net974),
    .S1(net987),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__mux4_1 clone7 (.A0(net804),
    .A1(net971),
    .A2(net1005),
    .A3(net789),
    .S0(net1013),
    .S1(net950),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net894),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net24),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net29),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net28),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_4 clone13 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net12),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_1 clone15 (.A(net11),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_1 clone16 (.A(net894),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net961),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net1046),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net998),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net998),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1039),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_1 clone22 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net29),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_1 clone27 (.A(net24),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net968),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1100),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_4 clone30 (.A(net921),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net7),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_1 clone32 (.A(net9),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net9),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_1 clone34 (.A(net6),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_1 clone35 (.A(net1087),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_1 clone36 (.A(net959),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_1 clone37 (.A(net997),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net959),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net1057),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net967),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net1104),
    .X(net1060));
 sky130_fd_sc_hd__buf_2 rebuffer42 (.A(clknet_1_0__leaf_net59),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net1061),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net526),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net535),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net540),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net651),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_1 fanout1 (.A(net969),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_1 fanout2 (.A(net932),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_1 fanout3 (.A(net971),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_1 fanout4 (.A(net977),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 fanout5 (.A(net987),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_1 fanout6 (.A(net1016),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_1 fanout7 (.A(net1013),
    .X(net1073));
 sky130_fd_sc_hd__buf_6 fanout8 (.A(net1005),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_1 fanout9 (.A(net985),
    .X(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in62));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in63));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(in64));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(in65));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(in66));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(in67));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(in68));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(in69));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(in70));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(in71));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(in72));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(in73));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(in74));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(in75));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(in76));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(in77));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(in78));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(in79));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(in80));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(in81));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(in82));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(in83));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(in84));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(in85));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(in86));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(in87));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(in88));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(in89));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(in90));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(in91));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(in92));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(in93));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(in94));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(in95));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(in96));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(in97));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(in98));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(in99));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A3 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_Q (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_S1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_Q_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_Q (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_X (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_S1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A0 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A3 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_S0 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_s824_D (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A3 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_Q_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_S0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_Q (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A3 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A3 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_S0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A0 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_X (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A3 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A2 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S0 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_s857_GATE (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A3 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_B1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_S0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A3 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A3 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_X (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_RESET_B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A4 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_X (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A3 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_X (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_Q (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_S0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A3 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_GATE (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_X (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A3 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net422_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge742_Q (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A3 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_S0 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A3 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A3 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A3 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_B1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_S1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge744_Q (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A2 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_A3 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A2 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_S0 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_Q (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S0 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_S1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge751_Q (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A3 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_X (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge752_Q_N (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge754_Q_N (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_s756_Q_N (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S0 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S0 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_s756_Q (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S0 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_s758_Q (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A3 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_S1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_S1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_s759_Q (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A2 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_S1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_s760_Q (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_S1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_S1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_S1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_s765_Q_N (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S0 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_S1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_S1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_s765_Q (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A3 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_S0 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_s766_Q (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_S1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_s768_Q (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A3 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_S0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_s770_Q (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A3 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_S0 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_s772_Q (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net544_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_s779_GCLK (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_s780_Q_N (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_S0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S0 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_s780_Q (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_S0 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_s783_Q (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_s784_Q (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_S0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_s785_Q (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A3 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S0 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_s787_Q (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A3 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_s788_Q (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A3 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_s789_Q_N (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_S1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_s789_Q (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_s792_Q (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A3 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_S1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_S1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_S1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_s796_Q_N (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A3 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A3 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_S1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_s796_Q (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A3 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A3 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_s799_Q (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A3 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_A3 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_s801_Q (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A3 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_S1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_S1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_S1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_S1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_s802_Q (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_S1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_S1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_s803_Q (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_s804_Q (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_s806_Q (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_S0 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A3 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_S0 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_S1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S0 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_S1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_S1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_s807_Q (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_S0 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S0 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_s812_Q_N (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_s819_Q (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_S0 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_S0 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_s828_Q_N (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S0 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_S1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_S0 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_S1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_s828_Q (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_S1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_S0 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_s831_Q (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S0 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_S1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_S1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_s832_Q (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_S1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A3 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_S1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_S1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_s833_Q (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A3 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S0 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A3 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_s834_Q (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_A3 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_S0 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_S1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_s835_Q (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_S1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_S0 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_s839_Q (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_S1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_S1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_S0 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_S1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_s840_Q (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_S0 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_s847_Q (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_s848_Q (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A3 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_S1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_s852_Q (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_S0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_s853_Q (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_S0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q_N (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_s860_Q (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_S0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_S1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_s863_Q (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A3 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_s869_Q (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A3 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_s880_Q (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c552_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_S1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_s887_Q (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_S0 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A2 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S0 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A3 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_S1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_s888_Q (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_S1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A3 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SET_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_A3 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_S1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_s892_Q (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S1 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_Q (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_S1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_Q_N (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A3 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_S1 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA_s928_Q (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_S0 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_Q (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_S0 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_S1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_Q (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_S0 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_S1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_Q (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S0 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_S1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_S1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_Q (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S0 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_S1 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A3 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_S1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_Q (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_S1 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_Q (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_S1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A4 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_RESET_B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A4 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A4 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_RESET_B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_RESET_B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_SCD (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_S0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_Q_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SCD (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_S1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_SCE (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_SCD (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A3 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_RESET_B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A3 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A3 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S0 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A3 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S0 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_X (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_S0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A3 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A0 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A0 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A2 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A2 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A0 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A0 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A3 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_S1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A3 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A2 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_S0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_S1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A2 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A0 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_A0 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_S1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A3 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A2 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A3 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c666_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A2 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S0 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A3 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A3 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_S0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A0 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A2 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_S0 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S0 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S0 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A3 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_S0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S0 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_X (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_X (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A3 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_X (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A2 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_X (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_X (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_X (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_A0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_X (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A2 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_X (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_A2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_X (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A3 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A2 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_X (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_X (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A3 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_X (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_S0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A0 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_X (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A1 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_X (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_S0 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_A1 (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_X (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_X (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_S1 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_X (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A3 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S1 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_X (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A3 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_S1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_A1 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_X (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_X (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A0 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_X (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A0 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A1 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_X (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S1 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A3 (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_X (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_s881_Q (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_S1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_S0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A1 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_A0 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A4 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_X (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_s775_Q (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A3 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_X (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_X (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_s836_Q (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_S1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net883_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_X (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_s781_Q (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_A2 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A3 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A1 (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_Q (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A1 (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_X (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_s798_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net908_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_s794_GCLK (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_S1 (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_c101_X (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_s808_Q (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S0 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_S0 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_X (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A2 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_S0 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A1 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_X (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A3 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_X (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_A (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A2 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_S0 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_A1 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_X (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_s771_Q (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_S1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S0 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A3 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A3 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A2 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A0 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_SCD (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A2 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A0 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A3 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A3 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCD (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c536_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A2 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A2 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_S0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_S1 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A0 (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_S0 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A3 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_S0 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A3 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A2 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A3 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A4 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A1 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_S0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_S0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A4 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_B1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_S0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_A0 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_S0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_SET_B (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A4 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A2 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A3 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A0 (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A1 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A2 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A3 (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer41_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_RESET_B (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_S0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c558_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A3 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_S0 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_S0 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_S0 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_S1 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_S1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer29_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer28_A (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A1 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S0 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A3 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A3 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S1 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_S1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_A3 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_S1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_S0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A2 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_S0 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_A2 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_S1 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_S0 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_S1 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A3 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A3 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_S1 (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_A1 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_S1 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_X (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c642_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S0 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A3 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S0 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A2 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_S0 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A1 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A4 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A3 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A4 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A3 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_S1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_S1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A3 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A4 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A4 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c640_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A0 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_A2 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A3 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S1 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S1 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_S0 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A3 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_S0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A2 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A4 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_S1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_S0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A3 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_B1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c128_A4 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_A0 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A2 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_X (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c527_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A3 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A0 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_S1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c116_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A4 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_S1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c638_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A3 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c264_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_B1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_s801_GATE_N (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s858_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s811_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s809_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s810_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s807_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s805_CLK (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s803_SLEEP_B (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_X (.DIODE(clknet_leaf_2_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s761_CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s826_CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_S0 (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_S1 (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S1 (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net888_X (.DIODE(clknet_1_0__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_S1 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_S0 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_S0 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_S0 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A2 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_S1 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A3 (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net888_X (.DIODE(clknet_1_1__leaf_net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_S1 (.DIODE(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A2 (.DIODE(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net618_X (.DIODE(clknet_1_1__leaf_net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A2 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A1 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net226_X (.DIODE(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A2 (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A3 (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A3 (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net226_X (.DIODE(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_S1 (.DIODE(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A3 (.DIODE(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A3 (.DIODE(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_S1 (.DIODE(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net596_X (.DIODE(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A1 (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A0 (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_A3 (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net204_X (.DIODE(clknet_1_0__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A2 (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_SET_B (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A1 (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A1 (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A0 (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A2 (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net204_X (.DIODE(clknet_1_1__leaf_net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A0 (.DIODE(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_A0 (.DIODE(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net411_X (.DIODE(clknet_1_1__leaf_net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net884_X (.DIODE(clknet_1_0__leaf_net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A3 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A0 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A0 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net142_X (.DIODE(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_A2 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A2 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A0 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A1 (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net142_X (.DIODE(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net342_X (.DIODE(clknet_1_1__leaf_net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net544_A (.DIODE(clknet_0_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net544_A (.DIODE(clknet_0_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net544_X (.DIODE(clknet_0_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_S1 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_S0 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A3 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net544_X (.DIODE(clknet_1_0__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_S1 (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_S1 (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SET_B (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A3 (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A1 (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net544_X (.DIODE(clknet_1_1__leaf_net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_B1 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A3 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A0 (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net291_X (.DIODE(clknet_1_0__leaf_net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_A2 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_A2 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A2 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A2 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A0 (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net299_X (.DIODE(clknet_1_0__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_SCD (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A1 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_S0 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A3 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S0 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A0 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A1 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_A2 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_c641_A0 (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net299_X (.DIODE(clknet_1_1__leaf_net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net883_A (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net883_A (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net883_X (.DIODE(clknet_0_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_A1 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S0 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SCD (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A2 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net883_X (.DIODE(clknet_1_0__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c281_S1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A2 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A0 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A2 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A3 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A2 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_S1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_S0 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A3 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_A3 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_A1 (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net883_X (.DIODE(clknet_1_1__leaf_net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A1 (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A3 (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A0 (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net114_X (.DIODE(clknet_1_1__leaf_net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net133_X (.DIODE(clknet_1_0__leaf_net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A2 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_A0 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A0 (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net899_X (.DIODE(clknet_1_1__leaf_net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_S1 (.DIODE(clknet_1_0__leaf_net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(clknet_1_0__leaf_net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(clknet_1_0__leaf_net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net115_X (.DIODE(clknet_1_0__leaf_net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A2 (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A1 (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A0 (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net207_X (.DIODE(clknet_1_1__leaf_net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net220_X (.DIODE(clknet_1_0__leaf_net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net897_A (.DIODE(clknet_0_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net897_A (.DIODE(clknet_0_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net897_X (.DIODE(clknet_0_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SCE (.DIODE(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A1 (.DIODE(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A3 (.DIODE(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net897_X (.DIODE(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A3 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A0 (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net897_X (.DIODE(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S1 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_S1 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_S1 (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net898_X (.DIODE(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A0 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S0 (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net898_X (.DIODE(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_S1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net62_X (.DIODE(clknet_1_0__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A3 (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A0 (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_S0 (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net62_X (.DIODE(clknet_1_1__leaf_net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer42_A (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A0 (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A2 (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A3 (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net59_X (.DIODE(clknet_1_0__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A0 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A3 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A0 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net59_X (.DIODE(clknet_1_1__leaf_net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_S0 (.DIODE(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A0 (.DIODE(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net57_X (.DIODE(clknet_1_0__leaf_net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_S1 (.DIODE(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_S0 (.DIODE(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net528_X (.DIODE(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_S1 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_S1 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_S1 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_S0 (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net528_X (.DIODE(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net47_A (.DIODE(clknet_0_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net47_A (.DIODE(clknet_0_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net47_X (.DIODE(clknet_0_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_S0 (.DIODE(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S1 (.DIODE(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_A0 (.DIODE(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net47_X (.DIODE(clknet_1_0__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A2 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net47_X (.DIODE(clknet_1_1__leaf_net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net882_A (.DIODE(clknet_0_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net882_A (.DIODE(clknet_0_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net882_X (.DIODE(clknet_0_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A1 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net882_X (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_A3 (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A1 (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_A0 (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net882_X (.DIODE(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_S0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A0 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone7_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_S0 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_X (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_S1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_SET_B (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_A0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_S0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer21_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone22_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer23_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A0 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_S0 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone27_X (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_X (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone34_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_D (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone35_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_S0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone5_A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A4 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_A0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_B1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_S0 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_S0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_SCE (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_A2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_S1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A3 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A3 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A0 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A0 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_X (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A3 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A0 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A3 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A3 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_A2 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_S1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_S1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_S0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_S0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_S0 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c530_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone4_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone3_A0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_S0 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_B1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_S0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_D (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_A0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_S1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_S0 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A3 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_X (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_X (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_SCE (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A0 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_X (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_S1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A3 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A0 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net1036));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net792),
    .A1(net789),
    .A2(net1009),
    .A3(net1084),
    .S0(net1069),
    .S1(net784),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net67),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1077),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net1078),
    .X(net1079));
 sky130_fd_sc_hd__mux4_1 clone6 (.A0(net1067),
    .A1(net25),
    .A2(net966),
    .A3(net1068),
    .S0(net1070),
    .S1(net1075),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net23),
    .X(net1081));
 sky130_fd_sc_hd__mux4_1 clone8 (.A0(net976),
    .A1(net964),
    .A2(net996),
    .A3(net965),
    .S0(net1101),
    .S1(net1071),
    .X(net1082));
 sky130_fd_sc_hd__mux4_1 clone9 (.A0(net804),
    .A1(net1069),
    .A2(net1074),
    .A3(net789),
    .S0(net1073),
    .S1(net950),
    .X(net1083));
 sky130_fd_sc_hd__mux4_1 clone10 (.A0(net958),
    .A1(net15),
    .A2(net1000),
    .A3(net990),
    .S0(net976),
    .S1(net978),
    .X(net1084));
 sky130_fd_sc_hd__a41o_1 clone11 (.A1(net5),
    .A2(net792),
    .A3(net778),
    .A4(net1002),
    .B1(net983),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net4),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net4),
    .X(net1087));
 sky130_fd_sc_hd__a41o_1 clone17 (.A1(net1101),
    .A2(net1075),
    .A3(net979),
    .A4(net990),
    .B1(net975),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_1 clone18 (.A(net894),
    .X(net1089));
 sky130_fd_sc_hd__a41o_1 clone19 (.A1(net978),
    .A2(net990),
    .A3(net979),
    .A4(net983),
    .B1(net1002),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(net12),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(net10),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_1 clone23 (.A(net16),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_1 clone24 (.A(net29),
    .X(net1094));
 sky130_fd_sc_hd__a41o_1 clone25 (.A1(net1072),
    .A2(net1018),
    .A3(net978),
    .A4(net983),
    .B1(net976),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(net8),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_1 clone28 (.A(net998),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 clone29 (.A(net847),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_1 clone33 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net10),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_1 clone39 (.A(net8),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_1 clone41 (.A(clknet_0_net62),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_1 clone42 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_1 clone43 (.A(net16),
    .X(net1104));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
