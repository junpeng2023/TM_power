module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net944;
 wire clknet_1_0__leaf_net944;
 wire clknet_1_1__leaf_net944;
 wire clknet_0_net696;
 wire clknet_1_0__leaf_net696;
 wire clknet_1_1__leaf_net696;
 wire clknet_0_net709;
 wire clknet_1_0__leaf_net709;
 wire clknet_1_1__leaf_net709;
 wire clknet_0_net858;
 wire clknet_1_0__leaf_net858;
 wire clknet_1_1__leaf_net858;
 wire clknet_0_net597;
 wire clknet_1_0__leaf_net597;
 wire clknet_1_1__leaf_net597;
 wire clknet_0_net611;
 wire clknet_1_0__leaf_net611;
 wire clknet_1_1__leaf_net611;
 wire clknet_0_net822;
 wire clknet_1_0__leaf_net822;
 wire clknet_1_1__leaf_net822;
 wire clknet_0_net994;
 wire clknet_1_0__leaf_net994;
 wire clknet_1_1__leaf_net994;
 wire clknet_0_net595;
 wire clknet_1_0__leaf_net595;
 wire clknet_1_1__leaf_net595;
 wire clknet_0_net607;
 wire clknet_1_0__leaf_net607;
 wire clknet_1_1__leaf_net607;
 wire clknet_0_net943;
 wire clknet_1_0__leaf_net943;
 wire clknet_1_1__leaf_net943;
 wire clknet_0_net703;
 wire clknet_1_0__leaf_net703;
 wire clknet_1_1__leaf_net703;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net942;
 wire clknet_1_0__leaf_net942;
 wire clknet_1_1__leaf_net942;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net570;
 wire clknet_1_0__leaf_net570;
 wire clknet_1_1__leaf_net570;
 wire clknet_0_net923;
 wire clknet_1_0__leaf_net923;
 wire clknet_1_1__leaf_net923;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net903;
 wire clknet_1_0__leaf_net903;
 wire clknet_1_1__leaf_net903;
 wire clknet_0_net902;
 wire clknet_1_0__leaf_net902;
 wire clknet_1_1__leaf_net902;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net596;
 wire clknet_1_0__leaf_net596;
 wire clknet_1_1__leaf_net596;
 wire clknet_0_net706;
 wire clknet_1_0__leaf_net706;
 wire clknet_1_1__leaf_net706;
 wire clknet_0_net562;
 wire clknet_1_0__leaf_net562;
 wire clknet_1_1__leaf_net562;
 wire clknet_0_net567;
 wire clknet_1_0__leaf_net567;
 wire clknet_1_1__leaf_net567;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net693;
 wire clknet_1_0__leaf_net693;
 wire clknet_1_1__leaf_net693;
 wire clknet_0_net561;
 wire clknet_1_0__leaf_net561;
 wire clknet_1_1__leaf_net561;
 wire clknet_0_net882;
 wire clknet_1_0__leaf_net882;
 wire clknet_1_1__leaf_net882;
 wire clknet_0_net700;
 wire clknet_1_0__leaf_net700;
 wire clknet_1_1__leaf_net700;
 wire clknet_0_net859;
 wire clknet_1_0__leaf_net859;
 wire clknet_1_1__leaf_net859;
 wire clknet_0_net436;
 wire clknet_1_0__leaf_net436;
 wire clknet_1_1__leaf_net436;
 wire clknet_0_net327;
 wire clknet_1_0__leaf_net327;
 wire clknet_1_1__leaf_net327;
 wire clknet_0_net313;
 wire clknet_1_0__leaf_net313;
 wire clknet_1_1__leaf_net313;
 wire clknet_0_net297;
 wire clknet_1_0__leaf_net297;
 wire clknet_1_1__leaf_net297;
 wire clknet_0_net881;
 wire clknet_1_0__leaf_net881;
 wire clknet_1_1__leaf_net881;
 wire clknet_0_net455;
 wire clknet_1_0__leaf_net455;
 wire clknet_1_1__leaf_net455;
 wire clknet_0_net985;
 wire clknet_1_0__leaf_net985;
 wire clknet_1_1__leaf_net985;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net286;
 wire clknet_1_0__leaf_net286;
 wire clknet_1_1__leaf_net286;
 wire clknet_0_net880;
 wire clknet_1_0__leaf_net880;
 wire clknet_1_1__leaf_net880;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net339;
 wire clknet_1_0__leaf_net339;
 wire clknet_1_1__leaf_net339;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net296;
 wire clknet_1_0__leaf_net296;
 wire clknet_1_1__leaf_net296;
 wire clknet_0_net823;
 wire clknet_1_0__leaf_net823;
 wire clknet_1_1__leaf_net823;
 wire clknet_0_net234;
 wire clknet_1_0__leaf_net234;
 wire clknet_1_1__leaf_net234;
 wire clknet_0_net225;
 wire clknet_1_0__leaf_net225;
 wire clknet_1_1__leaf_net225;
 wire clknet_0_net222;
 wire clknet_1_0__leaf_net222;
 wire clknet_1_1__leaf_net222;
 wire clknet_0_net499;
 wire clknet_1_0__leaf_net499;
 wire clknet_1_1__leaf_net499;
 wire clknet_0_net231;
 wire clknet_1_0__leaf_net231;
 wire clknet_1_1__leaf_net231;
 wire clknet_0_net226;
 wire clknet_1_0__leaf_net226;
 wire clknet_1_1__leaf_net226;
 wire clknet_0_net233;
 wire clknet_1_0__leaf_net233;
 wire clknet_1_1__leaf_net233;
 wire clknet_0_net819;
 wire clknet_1_0__leaf_net819;
 wire clknet_1_1__leaf_net819;
 wire clknet_0_net331;
 wire clknet_1_0__leaf_net331;
 wire clknet_1_1__leaf_net331;
 wire clknet_0_net635;
 wire clknet_1_0__leaf_net635;
 wire clknet_1_1__leaf_net635;
 wire clknet_0_net996;
 wire clknet_1_0__leaf_net996;
 wire clknet_1_1__leaf_net996;
 wire clknet_0_net352;
 wire clknet_1_0__leaf_net352;
 wire clknet_1_1__leaf_net352;
 wire clknet_0_net496;
 wire clknet_1_0__leaf_net496;
 wire clknet_1_1__leaf_net496;
 wire clknet_0_net309;
 wire clknet_1_0__leaf_net309;
 wire clknet_1_1__leaf_net309;
 wire clknet_0_net289;
 wire clknet_1_0__leaf_net289;
 wire clknet_1_1__leaf_net289;
 wire clknet_0_net489;
 wire clknet_1_0__leaf_net489;
 wire clknet_1_1__leaf_net489;
 wire clknet_0_net609;
 wire clknet_1_0__leaf_net609;
 wire clknet_1_1__leaf_net609;
 wire clknet_0_net605;
 wire clknet_1_0__leaf_net605;
 wire clknet_1_1__leaf_net605;
 wire clknet_0_net604;
 wire clknet_1_0__leaf_net604;
 wire clknet_1_1__leaf_net604;
 wire clknet_0_net470;
 wire clknet_1_0__leaf_net470;
 wire clknet_1_1__leaf_net470;
 wire clknet_0_net500;
 wire clknet_1_0__leaf_net500;
 wire clknet_1_1__leaf_net500;
 wire clknet_0_net504;
 wire clknet_1_0__leaf_net504;
 wire clknet_1_1__leaf_net504;
 wire clknet_0_net469;
 wire clknet_1_0__leaf_net469;
 wire clknet_1_1__leaf_net469;
 wire clknet_0_net442;
 wire clknet_1_0__leaf_net442;
 wire clknet_1_1__leaf_net442;
 wire clknet_0_net447;
 wire clknet_1_0__leaf_net447;
 wire clknet_1_1__leaf_net447;
 wire clknet_0_net163;
 wire clknet_1_0__leaf_net163;
 wire clknet_1_1__leaf_net163;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net317;
 wire clknet_1_0__leaf_net317;
 wire clknet_1_1__leaf_net317;
 wire clknet_0_net315;
 wire clknet_1_0__leaf_net315;
 wire clknet_1_1__leaf_net315;
 wire clknet_0_net221;
 wire clknet_1_0__leaf_net221;
 wire clknet_1_1__leaf_net221;
 wire clknet_0_net192;
 wire clknet_1_0__leaf_net192;
 wire clknet_1_1__leaf_net192;
 wire clknet_0_net174;
 wire clknet_1_0__leaf_net174;
 wire clknet_1_1__leaf_net174;
 wire clknet_0_net456;
 wire clknet_1_0__leaf_net456;
 wire clknet_1_1__leaf_net456;
 wire clknet_0_net320;
 wire clknet_1_0__leaf_net320;
 wire clknet_1_1__leaf_net320;
 wire clknet_0_net186;
 wire clknet_1_0__leaf_net186;
 wire clknet_1_1__leaf_net186;
 wire clknet_0_net185;
 wire clknet_1_0__leaf_net185;
 wire clknet_1_1__leaf_net185;
 wire clknet_0_net181;
 wire clknet_1_0__leaf_net181;
 wire clknet_1_1__leaf_net181;
 wire clknet_0_net175;
 wire clknet_1_0__leaf_net175;
 wire clknet_1_1__leaf_net175;
 wire clknet_0_net152;
 wire clknet_1_0__leaf_net152;
 wire clknet_1_1__leaf_net152;
 wire clknet_0_net167;
 wire clknet_1_0__leaf_net167;
 wire clknet_1_1__leaf_net167;
 wire clknet_0_net177;
 wire clknet_1_0__leaf_net177;
 wire clknet_1_1__leaf_net177;
 wire clknet_0_net600;
 wire clknet_1_0__leaf_net600;
 wire clknet_1_1__leaf_net600;
 wire clknet_0_net351;
 wire clknet_1_0__leaf_net351;
 wire clknet_1_1__leaf_net351;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net182;
 wire clknet_1_0__leaf_net182;
 wire clknet_1_1__leaf_net182;
 wire clknet_0_net179;
 wire clknet_1_0__leaf_net179;
 wire clknet_1_1__leaf_net179;
 wire clknet_0_net165;
 wire clknet_1_0__leaf_net165;
 wire clknet_1_1__leaf_net165;
 wire clknet_0_net191;
 wire clknet_1_0__leaf_net191;
 wire clknet_1_1__leaf_net191;
 wire clknet_0_net203;
 wire clknet_1_0__leaf_net203;
 wire clknet_1_1__leaf_net203;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net161;
 wire clknet_1_0__leaf_net161;
 wire clknet_1_1__leaf_net161;
 wire clknet_0_net437;
 wire clknet_1_0__leaf_net437;
 wire clknet_1_1__leaf_net437;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;

 sky130_fd_sc_hd__a31o_2 c100 (.A1(net30),
    .A2(net53),
    .A3(net62),
    .B1(net1034),
    .X(net70));
 sky130_fd_sc_hd__a21bo_1 c101 (.A1(net65),
    .A2(net63),
    .B1_N(net69),
    .X(net71));
 sky130_fd_sc_hd__a21bo_1 c102 (.A1(net1047),
    .A2(net65),
    .B1_N(net62),
    .X(net72));
 sky130_fd_sc_hd__xnor2_1 c103 (.A(net44),
    .B(net70),
    .Y(net73));
 sky130_fd_sc_hd__a21bo_1 c104 (.A1(net53),
    .A2(net1001),
    .B1_N(net71),
    .X(net74));
 sky130_fd_sc_hd__a21bo_1 c105 (.A1(net73),
    .A2(net47),
    .B1_N(net1034),
    .X(net75));
 sky130_fd_sc_hd__a21bo_4 c106 (.A1(net75),
    .A2(net62),
    .B1_N(net61),
    .X(net76));
 sky130_fd_sc_hd__a21bo_4 c107 (.A1(net1072),
    .A2(net74),
    .B1_N(net64),
    .X(net77));
 sky130_fd_sc_hd__mux4_2 c108 (.A0(net71),
    .A1(net1062),
    .A2(net76),
    .A3(net77),
    .S0(net23),
    .S1(net73),
    .X(net78));
 sky130_fd_sc_hd__xnor2_1 c109 (.A(net78),
    .B(net29),
    .Y(net79));
 sky130_fd_sc_hd__a21bo_1 c110 (.A1(net1060),
    .A2(net1052),
    .B1_N(net75),
    .X(net80));
 sky130_fd_sc_hd__xnor2_1 c111 (.A(net68),
    .B(net67),
    .Y(net81));
 sky130_fd_sc_hd__a41o_4 c112 (.A1(net1144),
    .A2(net63),
    .A3(net29),
    .A4(net70),
    .B1(net1029),
    .X(net82));
 sky130_fd_sc_hd__xnor2_1 c113 (.A(net64),
    .B(net1029),
    .Y(net83));
 sky130_fd_sc_hd__xnor2_4 c114 (.A(net76),
    .B(net77),
    .Y(net84));
 sky130_fd_sc_hd__a21bo_1 c115 (.A1(net75),
    .A2(net32),
    .B1_N(net19),
    .X(net85));
 sky130_fd_sc_hd__xnor2_1 c116 (.A(net80),
    .B(net84),
    .Y(net86));
 sky130_fd_sc_hd__xnor2_1 c117 (.A(net56),
    .B(net82),
    .Y(net87));
 sky130_fd_sc_hd__xnor2_4 c118 (.A(net1082),
    .B(net1021),
    .Y(net88));
 sky130_fd_sc_hd__a41o_1 c119 (.A1(net1091),
    .A2(net1029),
    .A3(net84),
    .A4(net72),
    .B1(net993),
    .X(net89));
 sky130_fd_sc_hd__a21bo_1 c120 (.A1(net29),
    .A2(net1037),
    .B1_N(net1101),
    .X(net90));
 sky130_fd_sc_hd__a21bo_1 c121 (.A1(net46),
    .A2(net67),
    .B1_N(net87),
    .X(net91));
 sky130_fd_sc_hd__a21bo_1 c122 (.A1(net1088),
    .A2(net89),
    .B1_N(net86),
    .X(net92));
 sky130_fd_sc_hd__a41o_1 c123 (.A1(net964),
    .A2(net87),
    .A3(net84),
    .A4(net68),
    .B1(net1029),
    .X(net93));
 sky130_fd_sc_hd__xnor2_1 c124 (.A(net93),
    .B(net1029),
    .Y(net94));
 sky130_fd_sc_hd__a41o_1 c125 (.A1(net89),
    .A2(net1060),
    .A3(net88),
    .A4(net93),
    .B1(net1029),
    .X(net95));
 sky130_fd_sc_hd__a41o_1 c126 (.A1(net32),
    .A2(net46),
    .A3(net1029),
    .A4(net88),
    .B1(net80),
    .X(net96));
 sky130_fd_sc_hd__a21bo_1 c127 (.A1(net87),
    .A2(net88),
    .B1_N(net90),
    .X(net97));
 sky130_fd_sc_hd__a21bo_1 c128 (.A1(net97),
    .A2(net84),
    .B1_N(net96),
    .X(net98));
 sky130_fd_sc_hd__a41o_2 c129 (.A1(net96),
    .A2(net94),
    .A3(net84),
    .A4(net1049),
    .B1(net75),
    .X(net99));
 sky130_fd_sc_hd__xnor2_4 c130 (.A(net99),
    .B(net82),
    .Y(net100));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net94),
    .A1(net98),
    .A2(net100),
    .A3(net86),
    .S0(net32),
    .S1(net99),
    .X(net101));
 sky130_fd_sc_hd__a21bo_2 c132 (.A1(net1105),
    .A2(net964),
    .B1_N(net1104),
    .X(net102));
 sky130_fd_sc_hd__a21bo_4 c133 (.A1(net1104),
    .A2(net1096),
    .B1_N(net1165),
    .X(net103));
 sky130_fd_sc_hd__xnor2_4 c134 (.A(net103),
    .B(net1097),
    .Y(net104));
 sky130_fd_sc_hd__xnor2_4 c135 (.A(net1095),
    .B(net1104),
    .Y(net105));
 sky130_fd_sc_hd__xnor2_4 c136 (.A(net1075),
    .B(net105),
    .Y(net106));
 sky130_fd_sc_hd__xnor2_4 c137 (.A(net968),
    .B(net1075),
    .Y(net107));
 sky130_fd_sc_hd__a21bo_4 c138 (.A1(net106),
    .A2(net1063),
    .B1_N(net1087),
    .X(net108));
 sky130_fd_sc_hd__a21bo_4 c139 (.A1(net108),
    .A2(net105),
    .B1_N(net1063),
    .X(net109));
 sky130_fd_sc_hd__a21bo_4 c140 (.A1(net968),
    .A2(net1054),
    .B1_N(net1104),
    .X(net110));
 sky130_fd_sc_hd__a31o_4 c141 (.A1(net110),
    .A2(net1063),
    .A3(net106),
    .B1(net1054),
    .X(net111));
 sky130_fd_sc_hd__a21bo_1 c142 (.A1(net1098),
    .A2(net1095),
    .B1_N(net111),
    .X(net112));
 sky130_fd_sc_hd__a21bo_4 c143 (.A1(net1044),
    .A2(net106),
    .B1_N(net1097),
    .X(net113));
 sky130_fd_sc_hd__a31o_4 c144 (.A1(net110),
    .A2(net113),
    .A3(net1044),
    .B1(net1063),
    .X(net114));
 sky130_fd_sc_hd__a21bo_1 c145 (.A1(net108),
    .A2(net110),
    .B1_N(net111),
    .X(net115));
 sky130_fd_sc_hd__a41o_4 c146 (.A1(net111),
    .A2(net1088),
    .A3(net110),
    .A4(net1044),
    .B1(net1094),
    .X(net116));
 sky130_fd_sc_hd__a31o_4 c147 (.A1(net114),
    .A2(net113),
    .A3(net1039),
    .B1(net1042),
    .X(net117));
 sky130_fd_sc_hd__a41o_4 c148 (.A1(net117),
    .A2(net1104),
    .A3(net103),
    .A4(net1039),
    .B1(net1042),
    .X(net118));
 sky130_fd_sc_hd__mux4_2 c149 (.A0(net117),
    .A1(net1044),
    .A2(net118),
    .A3(net106),
    .S0(net1102),
    .S1(net1100),
    .X(net119));
 sky130_fd_sc_hd__mux4_2 c150 (.A0(net118),
    .A1(net114),
    .A2(net113),
    .A3(net106),
    .S0(net1075),
    .S1(net1028),
    .X(net120));
 sky130_fd_sc_hd__mux4_2 c151 (.A0(net111),
    .A1(net120),
    .A2(net1044),
    .A3(net1091),
    .S0(net1102),
    .S1(net1028),
    .X(net121));
 sky130_fd_sc_hd__a31o_4 c152 (.A1(net120),
    .A2(net121),
    .A3(net1092),
    .B1(net1028),
    .X(net122));
 sky130_fd_sc_hd__mux4_2 c153 (.A0(net1028),
    .A1(net117),
    .A2(net120),
    .A3(net122),
    .S0(net105),
    .S1(net121),
    .X(net123));
 sky130_fd_sc_hd__a21bo_4 c154 (.A1(net114),
    .A2(net977),
    .B1_N(net979),
    .X(net124));
 sky130_fd_sc_hd__a21bo_2 c155 (.A1(net110),
    .A2(net1103),
    .B1_N(net1061),
    .X(net125));
 sky130_fd_sc_hd__a21bo_4 c156 (.A1(net1106),
    .A2(net103),
    .B1_N(net1102),
    .X(net126));
 sky130_fd_sc_hd__xnor2_4 c157 (.A(net118),
    .B(net979),
    .Y(net127));
 sky130_fd_sc_hd__a21bo_2 c158 (.A1(net113),
    .A2(net111),
    .B1_N(net1104),
    .X(net128));
 sky130_fd_sc_hd__a21bo_2 c159 (.A1(net127),
    .A2(net106),
    .B1_N(net1092),
    .X(net129));
 sky130_fd_sc_hd__mux4_2 c160 (.A0(net1107),
    .A1(net129),
    .A2(net126),
    .A3(net1028),
    .S0(net1147),
    .S1(net128),
    .X(net992));
 sky130_fd_sc_hd__a41o_4 c161 (.A1(net1097),
    .A2(net126),
    .A3(net124),
    .A4(net8),
    .B1(net1096),
    .X(net130));
 sky130_fd_sc_hd__xnor2_4 c162 (.A(net124),
    .B(net15),
    .Y(net131));
 sky130_fd_sc_hd__a21bo_2 c163 (.A1(net121),
    .A2(net129),
    .B1_N(net1165),
    .X(net132));
 sky130_fd_sc_hd__a21bo_4 c164 (.A1(net1106),
    .A2(net1082),
    .B1_N(net1089),
    .X(net133));
 sky130_fd_sc_hd__a21bo_4 c165 (.A1(net11),
    .A2(net133),
    .B1_N(net1027),
    .X(net134));
 sky130_fd_sc_hd__a41o_4 c166 (.A1(net108),
    .A2(net1173),
    .A3(net979),
    .A4(net129),
    .B1(net124),
    .X(net135));
 sky130_fd_sc_hd__xnor2_4 c167 (.A(net135),
    .B(net126),
    .Y(net136));
 sky130_fd_sc_hd__a21bo_4 c168 (.A1(net130),
    .A2(net132),
    .B1_N(net133),
    .X(net137));
 sky130_fd_sc_hd__a41o_2 c169 (.A1(net964),
    .A2(net137),
    .A3(net132),
    .A4(net1098),
    .B1(net126),
    .X(net138));
 sky130_fd_sc_hd__mux4_2 c170 (.A0(net129),
    .A1(net1130),
    .A2(net131),
    .A3(net1132),
    .S0(net130),
    .S1(net1073),
    .X(net139));
 sky130_fd_sc_hd__a41o_2 c171 (.A1(net1087),
    .A2(net132),
    .A3(net137),
    .A4(net1086),
    .B1(net1179),
    .X(net140));
 sky130_fd_sc_hd__a41o_4 c172 (.A1(net140),
    .A2(net128),
    .A3(net135),
    .A4(net15),
    .B1(net1086),
    .X(net141));
 sky130_fd_sc_hd__a41o_4 c173 (.A1(net1144),
    .A2(net134),
    .A3(net126),
    .A4(net1179),
    .B1(net131),
    .X(net142));
 sky130_fd_sc_hd__a41o_1 c174 (.A1(net137),
    .A2(net141),
    .A3(net140),
    .A4(net142),
    .B1(net138),
    .X(net143));
 sky130_fd_sc_hd__a41o_2 c175 (.A1(net141),
    .A2(net143),
    .A3(net140),
    .A4(net135),
    .B1(net1103),
    .X(net144));
 sky130_fd_sc_hd__xnor2_1 c176 (.A(net9),
    .B(net122),
    .Y(net145));
 sky130_fd_sc_hd__a31o_1 c177 (.A1(net144),
    .A2(net142),
    .A3(net132),
    .B1(net1020),
    .X(net146));
 sky130_fd_sc_hd__xnor2_2 c178 (.A(net1103),
    .B(net22),
    .Y(net147));
 sky130_fd_sc_hd__a31o_4 c179 (.A1(net1111),
    .A2(net1039),
    .A3(net1105),
    .B1(net1057),
    .X(net148));
 sky130_fd_sc_hd__a41o_4 c180 (.A1(net16),
    .A2(net114),
    .A3(net10),
    .A4(net0),
    .B1(net120),
    .X(net149));
 sky130_fd_sc_hd__a31o_2 c181 (.A1(net132),
    .A2(net141),
    .A3(net139),
    .B1(net1105),
    .X(net150));
 sky130_fd_sc_hd__mux4_2 c182 (.A0(net1052),
    .A1(net120),
    .A2(net1088),
    .A3(net977),
    .S0(net1057),
    .S1(net17),
    .X(net151));
 sky130_fd_sc_hd__a31o_1 c183 (.A1(net106),
    .A2(net1099),
    .A3(net149),
    .B1(clknet_1_1__leaf_net819),
    .X(net152));
 sky130_fd_sc_hd__xnor2_4 c184 (.A(net28),
    .B(net11),
    .Y(net153));
 sky130_fd_sc_hd__a21bo_1 c185 (.A1(net1165),
    .A2(net36),
    .B1_N(net1050),
    .X(net154));
 sky130_fd_sc_hd__a31o_2 c186 (.A1(net151),
    .A2(net145),
    .A3(net111),
    .B1(net1057),
    .X(net155));
 sky130_fd_sc_hd__a21bo_1 c187 (.A1(net1050),
    .A2(net124),
    .B1_N(net1057),
    .X(net156));
 sky130_fd_sc_hd__a41o_2 c188 (.A1(net154),
    .A2(net156),
    .A3(net1057),
    .A4(net1107),
    .B1(net1137),
    .X(net157));
 sky130_fd_sc_hd__a21bo_2 c189 (.A1(net1061),
    .A2(net154),
    .B1_N(net148),
    .X(net158));
 sky130_fd_sc_hd__a41o_4 c190 (.A1(net149),
    .A2(net1094),
    .A3(net157),
    .A4(net150),
    .B1(net124),
    .X(net159));
 sky130_fd_sc_hd__a21bo_1 c191 (.A1(net1045),
    .A2(net154),
    .B1_N(net1037),
    .X(net160));
 sky130_fd_sc_hd__a31o_1 c192 (.A1(clknet_1_1__leaf_net152),
    .A2(net20),
    .A3(net155),
    .B1(net1112),
    .X(net161));
 sky130_fd_sc_hd__mux4_2 c193 (.A0(net31),
    .A1(net28),
    .A2(net158),
    .A3(net135),
    .S0(net132),
    .S1(net1057),
    .X(net162));
 sky130_fd_sc_hd__a21bo_1 c194 (.A1(net17),
    .A2(net1050),
    .B1_N(clknet_1_1__leaf_net819),
    .X(net163));
 sky130_fd_sc_hd__a41o_2 c195 (.A1(net124),
    .A2(net156),
    .A3(net129),
    .A4(net1024),
    .B1(net162),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 c196 (.A0(net1024),
    .A1(net1097),
    .A2(net164),
    .A3(clknet_1_0__leaf_net152),
    .S0(net151),
    .S1(net162),
    .X(net165));
 sky130_fd_sc_hd__mux4_2 c197 (.A0(net145),
    .A1(net27),
    .A2(net21),
    .A3(net1057),
    .S0(net1045),
    .S1(net1024),
    .X(net166));
 sky130_fd_sc_hd__a41o_1 c198 (.A1(clknet_1_0__leaf_net152),
    .A2(net1089),
    .A3(net975),
    .A4(net31),
    .B1(net1054),
    .X(net167));
 sky130_fd_sc_hd__a41o_1 c199 (.A1(net1020),
    .A2(net27),
    .A3(net1137),
    .A4(net1031),
    .B1(net1102),
    .X(net168));
 sky130_fd_sc_hd__a41o_1 c200 (.A1(net992),
    .A2(net36),
    .A3(net51),
    .A4(net1089),
    .B1(net1048),
    .X(net169));
 sky130_fd_sc_hd__xnor2_1 c201 (.A(net156),
    .B(net51),
    .Y(net170));
 sky130_fd_sc_hd__xnor2_2 c202 (.A(net154),
    .B(net976),
    .Y(net171));
 sky130_fd_sc_hd__a31o_1 c203 (.A1(net102),
    .A2(net11),
    .A3(net1033),
    .B1(net1094),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 c204 (.A0(net1046),
    .A1(net1041),
    .A2(net43),
    .A3(net157),
    .S0(net168),
    .S1(net1020),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net145),
    .A1(net173),
    .A2(clknet_1_1__leaf_net163),
    .A3(net1031),
    .S0(net1049),
    .S1(net36),
    .X(net174));
 sky130_fd_sc_hd__a41o_1 c206 (.A1(net173),
    .A2(net1023),
    .A3(net1103),
    .A4(net172),
    .B1(clknet_1_0__leaf_net174),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 c207 (.A0(net151),
    .A1(net58),
    .A2(net54),
    .A3(net1046),
    .S0(net171),
    .S1(net1023),
    .X(net176));
 sky130_fd_sc_hd__a21bo_1 c208 (.A1(clknet_1_0__leaf_net167),
    .A2(net44),
    .B1_N(net1101),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 c209 (.A0(net176),
    .A1(net142),
    .A2(net1146),
    .A3(clknet_1_0__leaf_net177),
    .S0(net1023),
    .S1(net1175),
    .X(net178));
 sky130_fd_sc_hd__a31o_1 c210 (.A1(net43),
    .A2(net1175),
    .A3(clknet_1_0__leaf_net178),
    .B1(net1023),
    .X(net179));
 sky130_fd_sc_hd__a41o_1 c211 (.A1(net1175),
    .A2(clknet_1_1__leaf_net175),
    .A3(net128),
    .A4(net42),
    .B1(clknet_1_0__leaf_net178),
    .X(net180));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(clknet_1_0__leaf_net177),
    .A1(net135),
    .A2(net1024),
    .A3(clknet_1_0__leaf_net178),
    .S0(clknet_1_0__leaf_net174),
    .S1(clknet_1_1__leaf_net179),
    .X(net181));
 sky130_fd_sc_hd__a41o_1 c213 (.A1(net38),
    .A2(net176),
    .A3(clknet_1_0__leaf_net178),
    .A4(net975),
    .B1(net168),
    .X(net182));
 sky130_fd_sc_hd__sdfbbn_2 c214 (.CLK_N(clknet_4_1_0_clk),
    .D(net49),
    .RESET_B(net172),
    .SCD(net1023),
    .SCE(clknet_1_0__leaf_net181),
    .SET_B(net1089),
    .Q(net184),
    .Q_N(net183));
 sky130_fd_sc_hd__a41o_1 c215 (.A1(clknet_1_0__leaf_net174),
    .A2(net170),
    .A3(net1023),
    .A4(net183),
    .B1(net1091),
    .X(net185));
 sky130_fd_sc_hd__mux4_1 c216 (.A0(net1173),
    .A1(clknet_1_0__leaf_net178),
    .A2(net1023),
    .A3(clknet_1_0__leaf_net177),
    .S0(net29),
    .S1(clknet_1_0__leaf_net174),
    .X(net186));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_1__leaf_net186),
    .A1(net172),
    .A2(net176),
    .A3(clknet_1_0__leaf_net174),
    .S0(clknet_1_0__leaf_net178),
    .S1(net1050),
    .X(net187));
 sky130_fd_sc_hd__a41o_1 c218 (.A1(clknet_1_0__leaf_net178),
    .A2(net184),
    .A3(clknet_1_0__leaf_net186),
    .A4(clknet_1_0__leaf_net177),
    .B1(clknet_1_0__leaf_net181),
    .X(net188));
 sky130_fd_sc_hd__a41o_1 c219 (.A1(net134),
    .A2(clknet_1_0__leaf_net186),
    .A3(net159),
    .A4(clknet_1_1__leaf_net167),
    .B1(net826),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 c220 (.A0(net172),
    .A1(net1144),
    .A2(net42),
    .A3(net1041),
    .S0(net1034),
    .S1(net977),
    .X(net190));
 sky130_fd_sc_hd__a21bo_1 c221 (.A1(net36),
    .A2(clknet_1_0__leaf_net165),
    .B1_N(net1057),
    .X(net191));
 sky130_fd_sc_hd__a41o_1 c222 (.A1(clknet_1_0__leaf_net179),
    .A2(clknet_1_1__leaf_net163),
    .A3(net23),
    .A4(net11),
    .B1(net1092),
    .X(net192));
 sky130_fd_sc_hd__a41o_1 c223 (.A1(net1072),
    .A2(net1062),
    .A3(net1041),
    .A4(net74),
    .B1(net11),
    .X(net193));
 sky130_fd_sc_hd__a21bo_1 c224 (.A1(net70),
    .A2(net1023),
    .B1_N(net825),
    .X(net194));
 sky130_fd_sc_hd__a31o_1 c225 (.A1(net58),
    .A2(net48),
    .A3(net1027),
    .B1(net826),
    .X(net195));
 sky130_fd_sc_hd__sdfbbn_1 c226 (.CLK_N(clknet_4_1_0_clk),
    .D(net1113),
    .RESET_B(clknet_1_1__leaf_net192),
    .SCD(net164),
    .SCE(net1101),
    .SET_B(net1039),
    .Q(net197),
    .Q_N(net196));
 sky130_fd_sc_hd__a41o_4 c227 (.A1(net135),
    .A2(net77),
    .A3(net1023),
    .A4(net964),
    .B1(net137),
    .X(net198));
 sky130_fd_sc_hd__a41o_1 c228 (.A1(net69),
    .A2(clknet_1_0__leaf_net191),
    .A3(net38),
    .A4(net1034),
    .B1(net826),
    .X(net199));
 sky130_fd_sc_hd__a21bo_1 c229 (.A1(clknet_1_1__leaf_net191),
    .A2(net1026),
    .B1_N(net198),
    .X(net200));
 sky130_fd_sc_hd__sdfbbp_1 c230 (.CLK(clknet_4_1_0_clk),
    .D(net190),
    .RESET_B(net198),
    .SCD(net57),
    .SCE(clknet_1_1__leaf_net200),
    .SET_B(net79),
    .Q(net202),
    .Q_N(net201));
 sky130_fd_sc_hd__mux4_1 c231 (.A0(net195),
    .A1(net23),
    .A2(clknet_1_1__leaf_net191),
    .A3(net36),
    .S0(net76),
    .S1(net48),
    .X(net203));
 sky130_fd_sc_hd__a31o_1 c232 (.A1(net142),
    .A2(net164),
    .A3(net159),
    .B1(net1027),
    .X(net204));
 sky130_fd_sc_hd__sdfbbn_1 c233 (.CLK_N(clknet_4_1_0_clk),
    .D(net199),
    .RESET_B(clknet_1_0__leaf_net177),
    .SCD(clknet_1_0__leaf_net191),
    .SCE(net59),
    .SET_B(clknet_1_0__leaf_net179),
    .Q(net206),
    .Q_N(net205));
 sky130_fd_sc_hd__a41o_2 c234 (.A1(net42),
    .A2(net1186),
    .A3(net205),
    .A4(net198),
    .B1(net58),
    .X(net207));
 sky130_fd_sc_hd__a41o_1 c235 (.A1(net168),
    .A2(net207),
    .A3(net195),
    .A4(net1026),
    .B1(net787),
    .X(net208));
 sky130_fd_sc_hd__a41o_1 c236 (.A1(clknet_1_0__leaf_net175),
    .A2(clknet_1_0__leaf_net203),
    .A3(net206),
    .A4(net44),
    .B1(net1138),
    .X(net209));
 sky130_fd_sc_hd__mux4_2 c237 (.A0(net194),
    .A1(net1057),
    .A2(net195),
    .A3(net20),
    .S0(net48),
    .S1(net137),
    .X(net210));
 sky130_fd_sc_hd__a21bo_2 c238 (.A1(net195),
    .A2(net787),
    .B1_N(net825),
    .X(net1002));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net23),
    .A1(clknet_1_1__leaf_net185),
    .A2(net1041),
    .A3(net1052),
    .S0(net36),
    .S1(net787),
    .X(net211));
 sky130_fd_sc_hd__sdfrbp_2 c240 (.CLK(clknet_4_1_0_clk),
    .D(net208),
    .RESET_B(net206),
    .SCD(clknet_1_0__leaf_net175),
    .SCE(net30),
    .Q(net213),
    .Q_N(net212));
 sky130_fd_sc_hd__a41o_1 c241 (.A1(net193),
    .A2(net202),
    .A3(net212),
    .A4(net205),
    .B1(net787),
    .X(net214));
 sky130_fd_sc_hd__mux4_1 c242 (.A0(net1135),
    .A1(net41),
    .A2(net45),
    .A3(net979),
    .S0(net100),
    .S1(net1036),
    .X(net215));
 sky130_fd_sc_hd__mux4_1 c243 (.A0(net98),
    .A1(net1024),
    .A2(net100),
    .A3(net82),
    .S0(clknet_1_0__leaf_net192),
    .S1(net76),
    .X(net216));
 sky130_fd_sc_hd__mux4_2 c244 (.A0(net41),
    .A1(net979),
    .A2(net205),
    .A3(net54),
    .S0(net72),
    .S1(net1026),
    .X(net217));
 sky130_fd_sc_hd__mux4_1 c245 (.A0(clknet_1_1__leaf_net192),
    .A1(net1106),
    .A2(net1029),
    .A3(net183),
    .S0(net1135),
    .S1(net214),
    .X(net218));
 sky130_fd_sc_hd__mux4_1 c246 (.A0(net72),
    .A1(net95),
    .A2(net159),
    .A3(net1052),
    .S0(net1105),
    .S1(net1024),
    .X(net219));
 sky130_fd_sc_hd__mux4_1 c247 (.A0(net86),
    .A1(net60),
    .A2(net98),
    .A3(net95),
    .S0(net100),
    .S1(net873),
    .X(net220));
 sky130_fd_sc_hd__mux4_1 c248 (.A0(net83),
    .A1(net95),
    .A2(clknet_1_0__leaf_net163),
    .A3(net198),
    .S0(net72),
    .S1(net1098),
    .X(net221));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net23),
    .A1(net90),
    .A2(net210),
    .A3(net1030),
    .S0(clknet_1_1__leaf_net823),
    .S1(net825),
    .X(net222));
 sky130_fd_sc_hd__xnor2_4 c25 (.A(net976),
    .B(net977),
    .Y(net0));
 sky130_fd_sc_hd__mux4_1 c250 (.A0(net26),
    .A1(clknet_1_0__leaf_net200),
    .A2(net62),
    .A3(net1073),
    .S0(net207),
    .S1(net1136),
    .X(net223));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net214),
    .A1(net83),
    .A2(net1073),
    .A3(net1133),
    .S0(net198),
    .S1(net1139),
    .X(net224));
 sky130_fd_sc_hd__mux4_2 c252 (.A0(net82),
    .A1(net26),
    .A2(net964),
    .A3(net91),
    .S0(net794),
    .S1(net877),
    .X(net999));
 sky130_fd_sc_hd__mux4_1 c253 (.A0(net224),
    .A1(net67),
    .A2(clknet_1_0__leaf_net222),
    .A3(net1043),
    .S0(net1041),
    .S1(clknet_1_0__leaf_net823),
    .X(net225));
 sky130_fd_sc_hd__mux4_1 c254 (.A0(net67),
    .A1(clknet_1_0__leaf_net222),
    .A2(net183),
    .A3(net1092),
    .S0(net1144),
    .S1(net877),
    .X(net226));
 sky130_fd_sc_hd__mux4_1 c255 (.A0(clknet_1_0__leaf_net200),
    .A1(clknet_1_0__leaf_net226),
    .A2(net1029),
    .A3(clknet_1_0__leaf_net222),
    .S0(net999),
    .S1(net794),
    .X(net227));
 sky130_fd_sc_hd__mux4_2 c256 (.A0(net217),
    .A1(net91),
    .A2(net1073),
    .A3(net1030),
    .S0(net1037),
    .S1(net825),
    .X(net1004));
 sky130_fd_sc_hd__mux4_1 c257 (.A0(clknet_1_0__leaf_net192),
    .A1(clknet_1_0__leaf_net222),
    .A2(net1004),
    .A3(clknet_1_0__leaf_net226),
    .S0(net764),
    .S1(clknet_1_0__leaf_net823),
    .X(net228));
 sky130_fd_sc_hd__mux4_1 c258 (.A0(net62),
    .A1(net61),
    .A2(net1041),
    .A3(net70),
    .S0(net993),
    .S1(net857),
    .X(net229));
 sky130_fd_sc_hd__mux4_1 c259 (.A0(net86),
    .A1(net61),
    .A2(net201),
    .A3(net1004),
    .S0(net224),
    .S1(net764),
    .X(net230));
 sky130_fd_sc_hd__a31o_4 c26 (.A1(net1092),
    .A2(net1088),
    .A3(net0),
    .B1(net1094),
    .X(net1));
 sky130_fd_sc_hd__mux4_1 c260 (.A0(net70),
    .A1(net1098),
    .A2(clknet_1_0__leaf_net222),
    .A3(net59),
    .S0(net26),
    .S1(net965),
    .X(net231));
 sky130_fd_sc_hd__mux4_2 c261 (.A0(net1138),
    .A1(net41),
    .A2(net82),
    .A3(net1029),
    .S0(net1092),
    .S1(net877),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 c262 (.A0(net206),
    .A1(clknet_1_0__leaf_net226),
    .A2(net41),
    .A3(net1004),
    .S0(net85),
    .S1(net857),
    .X(net233));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net61),
    .A1(net85),
    .A2(net232),
    .A3(net1134),
    .S0(net1052),
    .S1(clknet_1_1__leaf_net823),
    .X(net234));
 sky130_fd_sc_hd__xnor2_4 c264 (.A(net1114),
    .B(net1132),
    .Y(net235));
 sky130_fd_sc_hd__xnor2_1 c265 (.A(net1091),
    .B(net103),
    .Y(net236));
 sky130_fd_sc_hd__xnor2_4 c266 (.A(net1042),
    .B(net118),
    .Y(net237));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net1142),
    .A2(net114),
    .B1_N(net1039),
    .X(net238));
 sky130_fd_sc_hd__a21bo_4 c268 (.A1(net1094),
    .A2(net1074),
    .B1_N(net1137),
    .X(net239));
 sky130_fd_sc_hd__xnor2_4 c269 (.A(net1074),
    .B(net235),
    .Y(net240));
 sky130_fd_sc_hd__xnor2_4 c27 (.A(net1),
    .B(net964),
    .Y(net2));
 sky130_fd_sc_hd__a21bo_4 c270 (.A1(net239),
    .A2(net103),
    .B1_N(net1137),
    .X(net241));
 sky130_fd_sc_hd__xnor2_4 c271 (.A(net241),
    .B(net1074),
    .Y(net242));
 sky130_fd_sc_hd__xnor2_4 c272 (.A(net122),
    .B(net1132),
    .Y(net243));
 sky130_fd_sc_hd__xnor2_4 c273 (.A(net1032),
    .B(net239),
    .Y(net244));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net240),
    .B(net244),
    .Y(net245));
 sky130_fd_sc_hd__mux4_2 c275 (.A0(net105),
    .A1(net241),
    .A2(net1074),
    .A3(net1092),
    .S0(net1032),
    .S1(net1015),
    .X(net246));
 sky130_fd_sc_hd__a21bo_4 c276 (.A1(net965),
    .A2(net243),
    .B1_N(net1032),
    .X(net247));
 sky130_fd_sc_hd__xnor2_4 c277 (.A(net244),
    .B(net243),
    .Y(net248));
 sky130_fd_sc_hd__a41o_4 c278 (.A1(net243),
    .A2(net244),
    .A3(net104),
    .A4(net1130),
    .B1(net1032),
    .X(net249));
 sky130_fd_sc_hd__a21bo_2 c279 (.A1(net239),
    .A2(net249),
    .B1_N(net248),
    .X(net250));
 sky130_fd_sc_hd__xnor2_4 c28 (.A(net968),
    .B(net1),
    .Y(net3));
 sky130_fd_sc_hd__mux4_1 c280 (.A0(net247),
    .A1(net1039),
    .A2(net240),
    .A3(net1012),
    .S0(net1032),
    .S1(net1102),
    .X(net251));
 sky130_fd_sc_hd__a41o_2 c281 (.A1(net241),
    .A2(net250),
    .A3(net1074),
    .A4(net244),
    .B1(net782),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 c282 (.A0(net1012),
    .A1(net252),
    .A2(net250),
    .A3(net237),
    .S0(net249),
    .X(net253));
 sky130_fd_sc_hd__a31o_4 c283 (.A1(net249),
    .A2(net252),
    .A3(net237),
    .B1(net783),
    .X(net254));
 sky130_fd_sc_hd__sdfbbn_2 c284 (.CLK_N(clknet_4_13_0_clk),
    .D(net248),
    .RESET_B(net1091),
    .SCD(net1012),
    .SCE(net1042),
    .SET_B(net783),
    .Q(net256),
    .Q_N(net255));
 sky130_fd_sc_hd__mux4_2 c285 (.A0(net250),
    .A1(net240),
    .A2(net256),
    .A3(net248),
    .S0(net235),
    .S1(net783),
    .X(net257));
 sky130_fd_sc_hd__xnor2_4 c286 (.A(net1015),
    .B(net1122),
    .Y(net258));
 sky130_fd_sc_hd__xnor2_4 c287 (.A(net1073),
    .B(net1086),
    .Y(net259));
 sky130_fd_sc_hd__a21bo_1 c288 (.A1(net1132),
    .A2(net968),
    .B1_N(net255),
    .X(net260));
 sky130_fd_sc_hd__xnor2_1 c289 (.A(net14),
    .B(net140),
    .Y(net261));
 sky130_fd_sc_hd__xnor2_4 c29 (.A(net979),
    .B(net975),
    .Y(net4));
 sky130_fd_sc_hd__a21bo_2 c290 (.A1(net15),
    .A2(net1087),
    .B1_N(net1018),
    .X(net262));
 sky130_fd_sc_hd__buf_2 c291 (.A(net1079),
    .X(net263));
 sky130_fd_sc_hd__a41o_1 c292 (.A1(net262),
    .A2(net1017),
    .A3(net144),
    .A4(net263),
    .B1(net119),
    .X(net264));
 sky130_fd_sc_hd__xnor2_2 c293 (.A(net1017),
    .B(net783),
    .Y(net265));
 sky130_fd_sc_hd__a21bo_1 c294 (.A1(net1042),
    .A2(net1017),
    .B1_N(net782),
    .X(net266));
 sky130_fd_sc_hd__a21bo_1 c295 (.A1(net266),
    .A2(net5),
    .B1_N(net1017),
    .X(net267));
 sky130_fd_sc_hd__xnor2_2 c296 (.A(net1184),
    .B(net250),
    .Y(net268));
 sky130_fd_sc_hd__mux4_2 c297 (.A0(net1102),
    .A1(net1103),
    .A2(net268),
    .A3(net143),
    .S0(net250),
    .S1(net1020),
    .X(net269));
 sky130_fd_sc_hd__a21bo_1 c298 (.A1(net248),
    .A2(net265),
    .B1_N(net1017),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 c299 (.A0(net126),
    .A1(net1017),
    .A2(net1010),
    .A3(net1015),
    .S0(net259),
    .S1(net3),
    .X(net271));
 sky130_fd_sc_hd__xnor2_1 c30 (.A(net975),
    .B(net968),
    .Y(net5));
 sky130_fd_sc_hd__xnor2_2 c300 (.A(net260),
    .B(net783),
    .Y(net272));
 sky130_fd_sc_hd__xnor2_2 c301 (.A(net252),
    .B(net272),
    .Y(net273));
 sky130_fd_sc_hd__a41o_1 c302 (.A1(net272),
    .A2(net2),
    .A3(net266),
    .A4(net1017),
    .B1(net241),
    .X(net274));
 sky130_fd_sc_hd__xnor2_1 c303 (.A(net143),
    .B(net257),
    .Y(net275));
 sky130_fd_sc_hd__mux4_1 c304 (.A0(net275),
    .A1(net274),
    .A2(net1015),
    .A3(net1184),
    .S0(net1010),
    .S1(net1153),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 c305 (.A0(net273),
    .A1(net244),
    .A2(net275),
    .A3(net1010),
    .S0(net1017),
    .S1(net6),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 c306 (.A0(net976),
    .A1(net144),
    .A2(net1010),
    .A3(net257),
    .S0(net828),
    .S1(net1078),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 c307 (.A0(net236),
    .A1(net138),
    .A2(net1012),
    .A3(net1010),
    .S0(net785),
    .S1(net1078),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 c308 (.A0(net1097),
    .A1(net149),
    .A2(net1094),
    .A3(net257),
    .S0(net1037),
    .S1(net1071),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 c309 (.A0(net267),
    .A1(net1097),
    .A2(net1035),
    .A3(net1129),
    .S0(net977),
    .S1(net1042),
    .X(net281));
 sky130_fd_sc_hd__xnor2_4 c31 (.A(net1084),
    .B(net968),
    .Y(net6));
 sky130_fd_sc_hd__mux4_1 c310 (.A0(net244),
    .A1(net254),
    .A2(net1183),
    .A3(net1102),
    .S0(net122),
    .S1(net785),
    .X(net282));
 sky130_fd_sc_hd__a41o_2 c311 (.A1(net129),
    .A2(net1018),
    .A3(net147),
    .A4(net1093),
    .B1(net1078),
    .X(net283));
 sky130_fd_sc_hd__sdfbbp_1 c312 (.CLK(clknet_4_4_0_clk),
    .D(net1183),
    .RESET_B(net269),
    .SCD(net255),
    .SCE(net258),
    .SET_B(clknet_1_1__leaf_net880),
    .Q(net285),
    .Q_N(net284));
 sky130_fd_sc_hd__a41o_1 c313 (.A1(net157),
    .A2(net1087),
    .A3(net1014),
    .A4(clknet_1_1__leaf_net859),
    .B1(clknet_1_0__leaf_net880),
    .X(net286));
 sky130_fd_sc_hd__sdfbbn_1 c314 (.CLK_N(clknet_4_12_0_clk),
    .D(net125),
    .RESET_B(net254),
    .SCD(net1050),
    .SCE(net283),
    .SET_B(net1078),
    .Q(net288),
    .Q_N(net287));
 sky130_fd_sc_hd__mux4_2 c315 (.A0(net128),
    .A1(net1020),
    .A2(net9),
    .A3(net1050),
    .S0(net1054),
    .S1(clknet_1_1__leaf_net819),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 c316 (.A0(net280),
    .A1(clknet_1_0__leaf_net286),
    .A2(net1131),
    .A3(net1010),
    .S0(net1038),
    .S1(net27),
    .X(net290));
 sky130_fd_sc_hd__sdfbbn_2 c317 (.CLK_N(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net286),
    .RESET_B(net243),
    .SCD(net109),
    .SCE(net267),
    .SET_B(net1014),
    .Q(net292),
    .Q_N(net291));
 sky130_fd_sc_hd__a41o_1 c318 (.A1(net1183),
    .A2(net111),
    .A3(net1099),
    .A4(net827),
    .B1(clknet_1_1__leaf_net880),
    .X(net293));
 sky130_fd_sc_hd__sdfbbp_1 c319 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net289),
    .RESET_B(net1010),
    .SCD(net157),
    .SCE(net1078),
    .SET_B(clknet_1_0__leaf_net880),
    .Q(net295),
    .Q_N(net294));
 sky130_fd_sc_hd__xnor2_4 c32 (.A(net1081),
    .B(net1),
    .Y(net7));
 sky130_fd_sc_hd__mux4_1 c320 (.A0(net1018),
    .A1(clknet_1_1__leaf_net293),
    .A2(net295),
    .A3(net284),
    .S0(net785),
    .S1(net1078),
    .X(net296));
 sky130_fd_sc_hd__mux4_1 c321 (.A0(clknet_1_0__leaf_net296),
    .A1(net127),
    .A2(clknet_1_1__leaf_net289),
    .A3(net147),
    .S0(clknet_1_0__leaf_net819),
    .S1(clknet_1_1__leaf_net859),
    .X(net297));
 sky130_fd_sc_hd__mux4_1 c322 (.A0(clknet_1_0__leaf_net161),
    .A1(net4),
    .A2(net147),
    .A3(net1020),
    .S0(net280),
    .S1(clknet_1_0__leaf_net880),
    .X(net298));
 sky130_fd_sc_hd__mux4_1 c323 (.A0(net254),
    .A1(clknet_1_0__leaf_net296),
    .A2(clknet_1_0__leaf_net297),
    .A3(clknet_1_1__leaf_net286),
    .S0(clknet_1_1__leaf_net293),
    .S1(net984),
    .X(net299));
 sky130_fd_sc_hd__mux4_1 c324 (.A0(clknet_1_1__leaf_net297),
    .A1(clknet_1_1__leaf_net293),
    .A2(net269),
    .A3(net1025),
    .S0(clknet_1_1__leaf_net286),
    .S1(clknet_1_1__leaf_net296),
    .X(net300));
 sky130_fd_sc_hd__a41o_1 c325 (.A1(clknet_1_0__leaf_net293),
    .A2(net128),
    .A3(net130),
    .A4(net294),
    .B1(clknet_1_1__leaf_net880),
    .X(net301));
 sky130_fd_sc_hd__mux4_1 c326 (.A0(net1071),
    .A1(clknet_1_1__leaf_net163),
    .A2(net1014),
    .A3(net259),
    .S0(net782),
    .S1(clknet_1_1__leaf_net881),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 c327 (.A0(net29),
    .A1(clknet_1_0__leaf_net302),
    .A2(net267),
    .A3(net239),
    .S0(net1015),
    .S1(clknet_1_0__leaf_net293),
    .X(net303));
 sky130_fd_sc_hd__a41o_1 c328 (.A1(net157),
    .A2(clknet_1_1__leaf_net302),
    .A3(net1014),
    .A4(net294),
    .B1(clknet_1_0__leaf_net882),
    .X(net304));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(clknet_1_0__leaf_net301),
    .A1(net159),
    .A2(clknet_1_1__leaf_net302),
    .A3(net842),
    .S0(clknet_1_1__leaf_net859),
    .S1(clknet_1_0__leaf_net882),
    .X(net305));
 sky130_fd_sc_hd__xnor2_2 c33 (.A(net964),
    .B(net968),
    .Y(net8));
 sky130_fd_sc_hd__mux4_1 c330 (.A0(net243),
    .A1(net57),
    .A2(net1055),
    .A3(net155),
    .S0(net1165),
    .S1(net24),
    .X(net306));
 sky130_fd_sc_hd__sdfbbn_2 c331 (.CLK_N(clknet_4_1_0_clk),
    .D(net144),
    .RESET_B(net166),
    .SCD(clknet_1_0__leaf_net178),
    .SCE(clknet_1_0__leaf_net302),
    .SET_B(clknet_1_0__leaf_net859),
    .Q(net308),
    .Q_N(net307));
 sky130_fd_sc_hd__mux4_1 c332 (.A0(net1131),
    .A1(net1091),
    .A2(net1031),
    .A3(net1018),
    .S0(net1014),
    .S1(clknet_1_1__leaf_net819),
    .X(net309));
 sky130_fd_sc_hd__a41o_1 c333 (.A1(net306),
    .A2(net292),
    .A3(net20),
    .A4(clknet_1_1__leaf_net163),
    .B1(net284),
    .X(net310));
 sky130_fd_sc_hd__sdfbbn_1 c334 (.CLK_N(clknet_4_6_0_clk),
    .D(net155),
    .RESET_B(net171),
    .SCD(net29),
    .SCE(clknet_1_0__leaf_net302),
    .SET_B(net1160),
    .Q(net312),
    .Q_N(net311));
 sky130_fd_sc_hd__a41o_1 c335 (.A1(clknet_1_1__leaf_net178),
    .A2(net1025),
    .A3(net243),
    .A4(net1137),
    .B1(clknet_1_0__leaf_net859),
    .X(net313));
 sky130_fd_sc_hd__mux4_1 c336 (.A0(clknet_1_1__leaf_net309),
    .A1(net295),
    .A2(net139),
    .A3(clknet_1_1__leaf_net313),
    .S0(net1095),
    .S1(clknet_1_0__leaf_net301),
    .X(net314));
 sky130_fd_sc_hd__a41o_1 c337 (.A1(net9),
    .A2(net51),
    .A3(clknet_1_1__leaf_net310),
    .A4(net291),
    .B1(net1023),
    .X(net315));
 sky130_fd_sc_hd__a41o_1 c338 (.A1(net170),
    .A2(net308),
    .A3(clknet_1_0__leaf_net301),
    .A4(clknet_1_0__leaf_net177),
    .B1(net785),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 c339 (.A0(net51),
    .A1(clknet_1_1__leaf_net310),
    .A2(net312),
    .A3(net294),
    .S0(net785),
    .S1(net1076),
    .X(net317));
 sky130_fd_sc_hd__a41o_4 c34 (.A1(net1081),
    .A2(net1060),
    .A3(net6),
    .A4(net1061),
    .B1(net1100),
    .X(net9));
 sky130_fd_sc_hd__mux4_1 c340 (.A0(clknet_1_0__leaf_net317),
    .A1(net311),
    .A2(net1039),
    .A3(clknet_1_1__leaf_net313),
    .S0(net141),
    .S1(net785),
    .X(net318));
 sky130_fd_sc_hd__mux4_1 c341 (.A0(net16),
    .A1(net257),
    .A2(clknet_1_1__leaf_net177),
    .A3(net38),
    .S0(clknet_1_1__leaf_net317),
    .S1(clknet_1_1__leaf_net178),
    .X(net319));
 sky130_fd_sc_hd__a41o_1 c342 (.A1(net1039),
    .A2(net292),
    .A3(net38),
    .A4(clknet_1_1__leaf_net174),
    .B1(net885),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 c343 (.A0(net148),
    .A1(clknet_1_0__leaf_net317),
    .A2(net307),
    .A3(net801),
    .S0(clknet_1_0__leaf_net819),
    .S1(net1076),
    .X(net321));
 sky130_fd_sc_hd__mux4_1 c344 (.A0(clknet_1_0__leaf_net317),
    .A1(clknet_1_0__leaf_net309),
    .A2(net965),
    .A3(clknet_1_0__leaf_net302),
    .S0(clknet_1_0__leaf_net177),
    .S1(net1027),
    .X(net322));
 sky130_fd_sc_hd__sdfbbp_1 c345 (.CLK(clknet_4_1_0_clk),
    .D(net312),
    .RESET_B(net1038),
    .SCD(clknet_1_1__leaf_net320),
    .SCE(clknet_1_0__leaf_net309),
    .SET_B(clknet_1_0__leaf_net819),
    .Q(net324),
    .Q_N(net323));
 sky130_fd_sc_hd__mux4_1 c346 (.A0(net128),
    .A1(net162),
    .A2(clknet_1_1__leaf_net320),
    .A3(net243),
    .S0(net984),
    .S1(net885),
    .X(net325));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net324),
    .A1(clknet_1_0__leaf_net309),
    .A2(net1048),
    .A3(net801),
    .S0(clknet_1_0__leaf_net859),
    .S1(net885),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c348 (.A0(net171),
    .A1(net311),
    .A2(net1185),
    .A3(net38),
    .S0(clknet_1_0__leaf_net174),
    .S1(clknet_1_0__leaf_net859),
    .X(net327));
 sky130_fd_sc_hd__a41o_1 c349 (.A1(clknet_1_0__leaf_net327),
    .A2(net306),
    .A3(clknet_1_1__leaf_net313),
    .A4(net885),
    .B1(net889),
    .X(net328));
 sky130_fd_sc_hd__xnor2_1 c35 (.A(net0),
    .B(net1081),
    .Y(net10));
 sky130_fd_sc_hd__mux4_1 c350 (.A0(clknet_1_1__leaf_net317),
    .A1(clknet_1_1__leaf_net327),
    .A2(net1019),
    .A3(net25),
    .S0(net801),
    .S1(net887),
    .X(net329));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net1035),
    .A1(clknet_1_0__leaf_net317),
    .A2(clknet_1_0__leaf_net309),
    .A3(clknet_1_0__leaf_net327),
    .S0(net801),
    .S1(net829),
    .X(net330));
 sky130_fd_sc_hd__a41o_1 c352 (.A1(net285),
    .A2(net1027),
    .A3(net78),
    .A4(net1082),
    .B1(clknet_1_0__leaf_net819),
    .X(net331));
 sky130_fd_sc_hd__mux4_1 c353 (.A0(clknet_1_0__leaf_net316),
    .A1(net1062),
    .A2(net1037),
    .A3(net1012),
    .S0(net1027),
    .S1(net826),
    .X(net332));
 sky130_fd_sc_hd__a41o_1 c354 (.A1(net207),
    .A2(net202),
    .A3(net148),
    .A4(net284),
    .B1(net307),
    .X(net333));
 sky130_fd_sc_hd__a21bo_1 c355 (.A1(net48),
    .A2(net292),
    .B1_N(net198),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 c356 (.A0(clknet_1_0__leaf_net310),
    .A1(net268),
    .A2(net1032),
    .A3(net210),
    .S0(net1088),
    .S1(net1024),
    .X(net335));
 sky130_fd_sc_hd__mux4_1 c357 (.A0(net169),
    .A1(clknet_1_1__leaf_net316),
    .A2(net1032),
    .A3(net1101),
    .S0(net183),
    .S1(net1043),
    .X(net336));
 sky130_fd_sc_hd__a31o_1 c358 (.A1(clknet_1_1__leaf_net181),
    .A2(net52),
    .A3(clknet_1_0__leaf_net313),
    .B1(net1047),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c359 (.A0(net52),
    .A1(net336),
    .A2(net268),
    .A3(net1138),
    .S0(net307),
    .S1(net988),
    .X(net338));
 sky130_fd_sc_hd__a21bo_4 c36 (.A1(net1072),
    .A2(net976),
    .B1_N(net1061),
    .X(net11));
 sky130_fd_sc_hd__mux4_1 c360 (.A0(net333),
    .A1(clknet_1_1__leaf_net174),
    .A2(net201),
    .A3(clknet_1_0__leaf_net316),
    .S0(net1054),
    .S1(net829),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c361 (.A0(net79),
    .A1(net308),
    .A2(net1024),
    .A3(clknet_1_0__leaf_net339),
    .S0(net52),
    .S1(net1022),
    .X(net340));
 sky130_fd_sc_hd__mux4_1 c362 (.A0(clknet_1_1__leaf_net316),
    .A1(net1148),
    .A2(net29),
    .A3(net1100),
    .S0(clknet_1_0__leaf_net310),
    .S1(net57),
    .X(net341));
 sky130_fd_sc_hd__mux4_1 c363 (.A0(net268),
    .A1(net24),
    .A2(net294),
    .A3(clknet_1_0__leaf_net339),
    .S0(net239),
    .S1(net891),
    .X(net342));
 sky130_fd_sc_hd__mux4_1 c364 (.A0(net57),
    .A1(net197),
    .A2(clknet_1_0__leaf_net339),
    .A3(clknet_1_1__leaf_net181),
    .S0(clknet_1_1__leaf_net177),
    .S1(net323),
    .X(net343));
 sky130_fd_sc_hd__a41o_1 c365 (.A1(net1057),
    .A2(clknet_1_1__leaf_net174),
    .A3(net1026),
    .A4(net872),
    .B1(net875),
    .X(net344));
 sky130_fd_sc_hd__sdfrbp_1 c366 (.CLK(clknet_4_3_0_clk),
    .D(net341),
    .RESET_B(net1152),
    .SCD(net166),
    .SCE(net1092),
    .Q(net346),
    .Q_N(net345));
 sky130_fd_sc_hd__mux4_1 c367 (.A0(net338),
    .A1(net1085),
    .A2(clknet_1_1__leaf_net174),
    .A3(clknet_1_0__leaf_net339),
    .S0(net54),
    .S1(net1024),
    .X(net347));
 sky130_fd_sc_hd__a41o_1 c368 (.A1(net335),
    .A2(net1052),
    .A3(net48),
    .A4(clknet_1_0__leaf_net339),
    .B1(net54),
    .X(net348));
 sky130_fd_sc_hd__a41o_1 c369 (.A1(net334),
    .A2(clknet_1_0__leaf_net339),
    .A3(net284),
    .A4(net164),
    .B1(net892),
    .X(net349));
 sky130_fd_sc_hd__xnor2_2 c37 (.A(net1100),
    .B(net1081),
    .Y(net12));
 sky130_fd_sc_hd__mux4_1 c370 (.A0(net30),
    .A1(net141),
    .A2(clknet_1_1__leaf_net181),
    .S0(net851),
    .S1(net892),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 c371 (.A0(clknet_1_1__leaf_net177),
    .A1(net295),
    .A2(net1101),
    .A3(net1039),
    .S0(net52),
    .S1(net792),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 c372 (.A0(clknet_1_1__leaf_net331),
    .A1(clknet_1_0__leaf_net351),
    .A2(net213),
    .A3(net1106),
    .S0(net792),
    .S1(net851),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net295),
    .A1(clknet_1_0__leaf_net165),
    .A2(net76),
    .A3(net1138),
    .S0(clknet_1_0__leaf_net339),
    .S1(clknet_1_1__leaf_net352),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 c374 (.A0(net45),
    .A1(net136),
    .A2(net91),
    .A3(net1099),
    .S0(net1034),
    .S1(net1026),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 c375 (.A0(net324),
    .A1(net1101),
    .A2(net88),
    .A3(clknet_1_0__leaf_net331),
    .S0(net198),
    .S1(net842),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 c376 (.A0(net20),
    .A1(net1024),
    .A2(net77),
    .A3(clknet_1_0__leaf_net185),
    .S0(net1089),
    .S1(net874),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 c377 (.A0(net37),
    .A1(clknet_1_0__leaf_net339),
    .A2(net60),
    .A3(net793),
    .S0(net842),
    .S1(net875),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 c378 (.A0(net37),
    .A1(net60),
    .A2(net1002),
    .A3(net1021),
    .S0(net77),
    .S1(net1106),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 c379 (.A0(net202),
    .A1(net90),
    .A2(net82),
    .A3(net1022),
    .S0(net210),
    .S1(net1089),
    .X(net359));
 sky130_fd_sc_hd__a21bo_4 c38 (.A1(net979),
    .A2(net4),
    .B1_N(net1083),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 c380 (.A0(net82),
    .A1(net45),
    .A2(clknet_1_0__leaf_net233),
    .A3(net1004),
    .S0(net88),
    .S1(net834),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 c381 (.A0(net82),
    .A1(net45),
    .A2(net1106),
    .A3(net88),
    .S0(net842),
    .S1(net857),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 c382 (.A0(net359),
    .A1(net358),
    .A2(clknet_1_0__leaf_net231),
    .A3(net130),
    .S0(clknet_1_0__leaf_net352),
    .S1(net1026),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 c383 (.A0(net230),
    .A1(net37),
    .A2(net229),
    .A3(net1026),
    .S0(net284),
    .S1(net1004),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 c384 (.A0(clknet_1_0__leaf_net185),
    .A1(clknet_1_1__leaf_net233),
    .A2(net90),
    .A3(net1026),
    .S0(net88),
    .S1(net765),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 c385 (.A0(net130),
    .A1(net92),
    .A2(net1103),
    .A3(net232),
    .S0(net857),
    .S1(clknet_1_0__leaf_net881),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 c386 (.A0(net85),
    .A1(net361),
    .A2(net285),
    .A3(clknet_1_1__leaf_net365),
    .S0(net999),
    .S1(clknet_1_0__leaf_net163),
    .X(net366));
 sky130_fd_sc_hd__mux4_1 c387 (.A0(net77),
    .A1(net37),
    .A2(clknet_1_1__leaf_net365),
    .A3(clknet_1_1__leaf_net185),
    .S0(clknet_1_0__leaf_net351),
    .S1(clknet_1_1__leaf_net366),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 c388 (.A0(clknet_1_1__leaf_net366),
    .A1(net20),
    .A2(net1101),
    .A3(net77),
    .S0(net1100),
    .S1(clknet_1_0__leaf_net881),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 c389 (.A0(net19),
    .A1(net1026),
    .A2(clknet_1_1__leaf_net366),
    .A3(net1052),
    .S0(clknet_1_1__leaf_net365),
    .S1(net1019),
    .X(net369));
 sky130_fd_sc_hd__xnor2_4 c39 (.A(net6),
    .B(net3),
    .Y(net14));
 sky130_fd_sc_hd__mux4_1 c390 (.A0(net363),
    .A1(clknet_1_0__leaf_net225),
    .A2(clknet_1_0__leaf_net365),
    .A3(net999),
    .S0(net834),
    .S1(net894),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 c391 (.A0(clknet_1_0__leaf_net163),
    .A1(net88),
    .A2(net1026),
    .A3(net323),
    .S0(clknet_1_1__leaf_net365),
    .S1(net893),
    .X(net371));
 sky130_fd_sc_hd__mux4_1 c392 (.A0(net91),
    .A1(net371),
    .A2(net230),
    .A3(clknet_1_0__leaf_net366),
    .S0(net100),
    .S1(net1019),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 c393 (.A0(net362),
    .A1(net1094),
    .A2(clknet_1_0__leaf_net366),
    .A3(clknet_1_0__leaf_net365),
    .S0(net808),
    .S1(net898),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 c394 (.A0(net54),
    .A1(net284),
    .A2(net45),
    .A3(net829),
    .S0(net893),
    .S1(net896),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 c395 (.A0(clknet_1_0__leaf_net365),
    .A1(clknet_1_0__leaf_net366),
    .A2(clknet_1_0__leaf_net352),
    .A3(net374),
    .S1(net897),
    .X(net375));
 sky130_fd_sc_hd__a41o_2 c396 (.A1(net1100),
    .A2(net1097),
    .A3(net1130),
    .A4(net1020),
    .B1(net1032),
    .X(net376));
 sky130_fd_sc_hd__xnor2_2 c397 (.A(net1108),
    .B(net249),
    .Y(net377));
 sky130_fd_sc_hd__xnor2_4 c398 (.A(net239),
    .B(net242),
    .Y(net378));
 sky130_fd_sc_hd__xnor2_2 c399 (.A(net1099),
    .B(net376),
    .Y(net379));
 sky130_fd_sc_hd__xnor2_4 c40 (.A(net7),
    .B(net1072),
    .Y(net15));
 sky130_fd_sc_hd__a21bo_2 c400 (.A1(net1140),
    .A2(net379),
    .B1_N(net1105),
    .X(net380));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net1098),
    .B(net256),
    .Y(net381));
 sky130_fd_sc_hd__xnor2_2 c402 (.A(net380),
    .B(net247),
    .Y(net382));
 sky130_fd_sc_hd__clkbuf_2 c403 (.A(net1079),
    .X(net383));
 sky130_fd_sc_hd__xnor2_2 c404 (.A(net1068),
    .B(net1016),
    .Y(net384));
 sky130_fd_sc_hd__a21bo_2 c405 (.A1(net1097),
    .A2(net383),
    .B1_N(net1067),
    .X(net385));
 sky130_fd_sc_hd__xnor2_1 c406 (.A(net1059),
    .B(net238),
    .Y(net386));
 sky130_fd_sc_hd__a21bo_2 c407 (.A1(net1120),
    .A2(net384),
    .B1_N(net1067),
    .X(net387));
 sky130_fd_sc_hd__mux4_2 c408 (.A0(net386),
    .A1(net107),
    .A2(net965),
    .A3(net109),
    .S0(net1059),
    .S1(net1068),
    .X(net388));
 sky130_fd_sc_hd__a31o_1 c409 (.A1(net1042),
    .A2(net386),
    .A3(net1059),
    .B1(net1067),
    .X(net389));
 sky130_fd_sc_hd__a41o_1 c41 (.A1(net1083),
    .A2(net15),
    .A3(net1056),
    .A4(net1097),
    .B1(net6),
    .X(net990));
 sky130_fd_sc_hd__mux4_2 c410 (.A0(net235),
    .A1(net1016),
    .A2(net380),
    .A3(net245),
    .S0(net1147),
    .S1(net1059),
    .X(net390));
 sky130_fd_sc_hd__a21bo_1 c411 (.A1(net389),
    .A2(net245),
    .B1_N(net1067),
    .X(net391));
 sky130_fd_sc_hd__a31o_1 c412 (.A1(net1016),
    .A2(net390),
    .A3(net247),
    .B1(net1059),
    .X(net392));
 sky130_fd_sc_hd__sdfbbn_2 c413 (.CLK_N(clknet_4_13_0_clk),
    .D(net122),
    .RESET_B(net387),
    .SCD(net1147),
    .SCE(net1067),
    .SET_B(net388),
    .Q(net394),
    .Q_N(net393));
 sky130_fd_sc_hd__mux4_2 c414 (.A0(net394),
    .A1(net377),
    .A2(net249),
    .A3(net380),
    .S0(net1068),
    .S1(net1042),
    .X(net395));
 sky130_fd_sc_hd__xnor2_4 c415 (.A(net394),
    .B(net766),
    .Y(net396));
 sky130_fd_sc_hd__a41o_1 c416 (.A1(net389),
    .A2(net388),
    .A3(net393),
    .A4(net1067),
    .B1(net1079),
    .X(net397));
 sky130_fd_sc_hd__a41o_2 c417 (.A1(net378),
    .A2(net377),
    .A3(net248),
    .A4(net383),
    .B1(net1079),
    .X(net398));
 sky130_fd_sc_hd__a41o_4 c418 (.A1(net266),
    .A2(net1140),
    .A3(net1147),
    .A4(net981),
    .B1(net1017),
    .X(net399));
 sky130_fd_sc_hd__a41o_4 c419 (.A1(net0),
    .A2(net266),
    .A3(net1147),
    .A4(net1067),
    .B1(net1076),
    .X(net400));
 sky130_fd_sc_hd__a41o_4 c42 (.A1(net1056),
    .A2(net1060),
    .A3(net15),
    .A4(net1052),
    .B1(net1093),
    .X(net16));
 sky130_fd_sc_hd__a31o_1 c420 (.A1(net1099),
    .A2(net379),
    .A3(net1018),
    .B1(net1078),
    .X(net401));
 sky130_fd_sc_hd__a41o_2 c421 (.A1(net265),
    .A2(net263),
    .A3(net239),
    .A4(net1018),
    .B1(net1079),
    .X(net402));
 sky130_fd_sc_hd__sdfbbn_2 c422 (.CLK_N(clknet_4_5_0_clk),
    .D(net250),
    .RESET_B(net241),
    .SCD(net1067),
    .SCE(net399),
    .SET_B(net252),
    .Q(net404),
    .Q_N(net403));
 sky130_fd_sc_hd__sdfrtn_1 c423 (.CLK_N(clknet_4_13_0_clk),
    .D(net275),
    .RESET_B(net378),
    .SCD(net138),
    .SCE(net1016),
    .Q(net405));
 sky130_fd_sc_hd__a41o_1 c424 (.A1(net1100),
    .A2(net1040),
    .A3(net1091),
    .A4(net403),
    .B1(net1076),
    .X(net406));
 sky130_fd_sc_hd__a21bo_1 c425 (.A1(net389),
    .A2(net138),
    .B1_N(net1045),
    .X(net407));
 sky130_fd_sc_hd__sdfrtp_4 c426 (.CLK(clknet_4_5_0_clk),
    .D(net399),
    .RESET_B(net272),
    .SCD(net274),
    .SCE(net400),
    .Q(net408));
 sky130_fd_sc_hd__a41o_1 c427 (.A1(net140),
    .A2(net400),
    .A3(net263),
    .A4(net403),
    .B1(net1042),
    .X(net409));
 sky130_fd_sc_hd__a41o_2 c428 (.A1(net241),
    .A2(net376),
    .A3(net1095),
    .A4(net1099),
    .B1(net827),
    .X(net410));
 sky130_fd_sc_hd__sdfbbp_1 c429 (.CLK(clknet_4_13_0_clk),
    .D(net139),
    .RESET_B(net406),
    .SCD(net133),
    .SCE(net387),
    .SET_B(net400),
    .Q(net412),
    .Q_N(net411));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net15),
    .A1(net9),
    .A2(net1056),
    .A3(net1052),
    .S0(net13),
    .S1(net1097),
    .X(net17));
 sky130_fd_sc_hd__sdfbbn_1 c430 (.CLK_N(clknet_4_5_0_clk),
    .D(net390),
    .RESET_B(net1080),
    .SCD(net391),
    .SCE(net269),
    .SET_B(net400),
    .Q(net414),
    .Q_N(net413));
 sky130_fd_sc_hd__a31o_1 c431 (.A1(net1080),
    .A2(net238),
    .A3(net265),
    .B1(net411),
    .X(net415));
 sky130_fd_sc_hd__a41o_1 c432 (.A1(net1130),
    .A2(net383),
    .A3(net1080),
    .A4(net403),
    .B1(net411),
    .X(net416));
 sky130_fd_sc_hd__sdfbbn_1 c433 (.CLK_N(clknet_4_12_0_clk),
    .D(net260),
    .RESET_B(net259),
    .SCD(net402),
    .SCE(net412),
    .SET_B(net1012),
    .Q(net418),
    .Q_N(net417));
 sky130_fd_sc_hd__a41o_1 c434 (.A1(net8),
    .A2(net410),
    .A3(net1127),
    .A4(net1080),
    .B1(net403),
    .X(net419));
 sky130_fd_sc_hd__a31o_2 c435 (.A1(net237),
    .A2(net416),
    .A3(net410),
    .B1(net1018),
    .X(net420));
 sky130_fd_sc_hd__mux4_1 c436 (.A0(net405),
    .A1(net237),
    .A2(net410),
    .A3(net1100),
    .S0(net415),
    .S1(net1080),
    .X(net421));
 sky130_fd_sc_hd__mux4_2 c437 (.A0(net401),
    .A1(net419),
    .A2(net412),
    .A3(net410),
    .S0(net403),
    .S1(net812),
    .X(net422));
 sky130_fd_sc_hd__mux4_1 c438 (.A0(net420),
    .A1(net241),
    .A2(net260),
    .A3(net414),
    .S0(net1080),
    .S1(net1008),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 c439 (.A0(net992),
    .A1(net419),
    .A2(net402),
    .A3(net265),
    .S0(net1008),
    .S1(net781),
    .X(net424));
 sky130_fd_sc_hd__xnor2_4 c44 (.A(net1101),
    .B(net1),
    .Y(net18));
 sky130_fd_sc_hd__mux4_1 c440 (.A0(net155),
    .A1(net254),
    .A2(net1008),
    .A3(net405),
    .S0(net1009),
    .S1(clknet_1_1__leaf_net881),
    .X(net425));
 sky130_fd_sc_hd__a21bo_1 c441 (.A1(net377),
    .A2(net125),
    .B1_N(net25),
    .X(net426));
 sky130_fd_sc_hd__a21bo_2 c442 (.A1(net977),
    .A2(net245),
    .B1_N(net854),
    .X(net427));
 sky130_fd_sc_hd__mux4_1 c443 (.A0(net269),
    .A1(net376),
    .A2(net1008),
    .A3(net1018),
    .S0(net263),
    .S1(net1161),
    .X(net428));
 sky130_fd_sc_hd__a21bo_1 c444 (.A1(net426),
    .A2(net1125),
    .B1_N(net812),
    .X(net429));
 sky130_fd_sc_hd__a31o_1 c445 (.A1(net376),
    .A2(net148),
    .A3(net410),
    .B1(net291),
    .X(net430));
 sky130_fd_sc_hd__a41o_1 c446 (.A1(net262),
    .A2(net1008),
    .A3(net1067),
    .A4(net798),
    .B1(net842),
    .X(net431));
 sky130_fd_sc_hd__a41o_1 c447 (.A1(net1080),
    .A2(net1086),
    .A3(net413),
    .A4(net1018),
    .B1(net854),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 c448 (.A0(net272),
    .A1(net416),
    .A2(net166),
    .A3(clknet_1_1__leaf_net165),
    .S0(net376),
    .S1(net1109),
    .X(net433));
 sky130_fd_sc_hd__mux4_2 c449 (.A0(net288),
    .A1(net150),
    .A2(net155),
    .A3(net1070),
    .S0(net1095),
    .S1(net781),
    .X(net434));
 sky130_fd_sc_hd__xnor2_1 c45 (.A(net1060),
    .B(net965),
    .Y(net19));
 sky130_fd_sc_hd__mux4_1 c450 (.A0(net433),
    .A1(clknet_1_0__leaf_net161),
    .A2(net1035),
    .A3(net422),
    .S0(net247),
    .S1(net1076),
    .X(net435));
 sky130_fd_sc_hd__a21bo_1 c451 (.A1(net398),
    .A2(clknet_1_1__leaf_net859),
    .B1_N(net1076),
    .X(net436));
 sky130_fd_sc_hd__a31o_1 c452 (.A1(net30),
    .A2(clknet_1_0__leaf_net161),
    .A3(net150),
    .B1(net854),
    .X(net437));
 sky130_fd_sc_hd__a21bo_1 c453 (.A1(net388),
    .A2(net1025),
    .B1_N(net780),
    .X(net438));
 sky130_fd_sc_hd__a41o_1 c454 (.A1(net416),
    .A2(clknet_1_1__leaf_net436),
    .A3(net403),
    .A4(net31),
    .B1(net410),
    .X(net439));
 sky130_fd_sc_hd__sdfbbp_1 c455 (.CLK(clknet_4_12_0_clk),
    .D(net109),
    .RESET_B(clknet_1_1__leaf_net437),
    .SCD(net438),
    .SCE(net434),
    .SET_B(net854),
    .Q(net441),
    .Q_N(net440));
 sky130_fd_sc_hd__mux4_1 c456 (.A0(net134),
    .A1(net438),
    .A2(net440),
    .A3(clknet_1_1__leaf_net289),
    .S0(net1096),
    .S1(net842),
    .X(net442));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net430),
    .A1(net259),
    .A2(clknet_1_0__leaf_net442),
    .A3(net24),
    .S0(net440),
    .S1(net899),
    .X(net443));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net443),
    .A1(net377),
    .A2(net259),
    .A3(clknet_1_0__leaf_net442),
    .S0(net440),
    .S1(net899),
    .X(net444));
 sky130_fd_sc_hd__mux4_1 c459 (.A0(net1080),
    .A1(clknet_1_1__leaf_net442),
    .A2(clknet_1_1__leaf_net436),
    .A3(net378),
    .S0(net799),
    .S1(net900),
    .X(net445));
 sky130_fd_sc_hd__xnor2_4 c46 (.A(net1103),
    .B(net1091),
    .Y(net20));
 sky130_fd_sc_hd__a41o_2 c460 (.A1(net138),
    .A2(net441),
    .A3(net799),
    .A4(net854),
    .B1(net900),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(clknet_1_1__leaf_net442),
    .A1(net138),
    .A2(net992),
    .A3(net446),
    .S0(net780),
    .S1(net854),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 c462 (.A0(net438),
    .A1(net14),
    .A2(net977),
    .A3(net1036),
    .S0(clknet_1_1__leaf_net177),
    .S1(net889),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 c463 (.A0(net1047),
    .A1(net1071),
    .A2(net402),
    .A3(clknet_1_1__leaf_net182),
    .S0(net1090),
    .S1(net900),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 c464 (.A0(net414),
    .A1(clknet_1_1__leaf_net317),
    .A2(net142),
    .A3(net1001),
    .S0(net1100),
    .S1(net886),
    .X(net450));
 sky130_fd_sc_hd__mux4_1 c465 (.A0(net308),
    .A1(clknet_1_1__leaf_net301),
    .A2(net1031),
    .A3(net434),
    .S0(net25),
    .S1(net890),
    .X(net451));
 sky130_fd_sc_hd__mux4_1 c466 (.A0(net27),
    .A1(net1048),
    .A2(net1141),
    .A3(net1091),
    .S0(clknet_1_1__leaf_net174),
    .S1(clknet_1_0__leaf_net902),
    .X(net452));
 sky130_fd_sc_hd__mux4_1 c467 (.A0(clknet_1_1__leaf_net313),
    .A1(net410),
    .A2(net393),
    .A3(net1053),
    .S0(net883),
    .S1(net889),
    .X(net453));
 sky130_fd_sc_hd__mux4_1 c468 (.A0(net429),
    .A1(clknet_1_0__leaf_net182),
    .A2(clknet_1_1__leaf_net302),
    .A3(net155),
    .S0(net403),
    .S1(net883),
    .X(net454));
 sky130_fd_sc_hd__mux4_1 c469 (.A0(net446),
    .A1(net1096),
    .A2(net413),
    .A3(net393),
    .S0(clknet_1_1__leaf_net881),
    .S1(net886),
    .X(net455));
 sky130_fd_sc_hd__xnor2_4 c47 (.A(net1051),
    .B(net1053),
    .Y(net21));
 sky130_fd_sc_hd__mux4_1 c470 (.A0(net1051),
    .A1(net977),
    .A2(net1001),
    .A3(net1185),
    .S0(net1031),
    .S1(clknet_1_0__leaf_net174),
    .X(net456));
 sky130_fd_sc_hd__mux4_1 c471 (.A0(net397),
    .A1(net245),
    .A2(net1093),
    .A3(net1038),
    .S0(clknet_1_1__leaf_net456),
    .S1(net866),
    .X(net457));
 sky130_fd_sc_hd__mux4_2 c472 (.A0(net1128),
    .A1(net245),
    .A2(net31),
    .A3(net50),
    .S0(net836),
    .S1(net884),
    .X(net458));
 sky130_fd_sc_hd__mux4_1 c473 (.A0(net256),
    .A1(net1014),
    .A2(clknet_1_1__leaf_net317),
    .A3(net410),
    .S0(net1106),
    .S1(clknet_1_0__leaf_net901),
    .X(net459));
 sky130_fd_sc_hd__mux4_1 c474 (.A0(net410),
    .A1(net397),
    .A2(net422),
    .A3(net1123),
    .S0(net27),
    .S1(net904),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 c475 (.A0(clknet_1_1__leaf_net302),
    .A1(net414),
    .A2(clknet_1_0__leaf_net436),
    .A3(net889),
    .S0(net890),
    .S1(net904),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 c476 (.A0(net134),
    .A1(net400),
    .A2(net399),
    .A3(net27),
    .S0(net835),
    .S1(net907),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 c477 (.A0(net397),
    .A1(net1098),
    .A2(net136),
    .A3(net1031),
    .S0(net835),
    .S1(net905),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net448),
    .A1(clknet_1_0__leaf_net182),
    .A2(clknet_1_1__leaf_net455),
    .A3(net900),
    .S0(net905),
    .S1(net908),
    .X(net985));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(clknet_1_0__leaf_net455),
    .A1(net1115),
    .A2(net16),
    .A3(net255),
    .S0(clknet_1_1__leaf_net985),
    .S1(net909),
    .X(net464));
 sky130_fd_sc_hd__xnor2_2 c48 (.A(net4),
    .B(net1173),
    .Y(net22));
 sky130_fd_sc_hd__mux4_2 c480 (.A0(net1025),
    .A1(net1094),
    .A2(net1036),
    .A3(net248),
    .S0(net803),
    .S1(net906),
    .X(net465));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net1032),
    .A1(net465),
    .A2(net142),
    .A3(net890),
    .S0(net900),
    .S1(net906),
    .X(net466));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_1__leaf_net182),
    .A1(clknet_1_0__leaf_net315),
    .A2(net466),
    .A3(clknet_1_0__leaf_net436),
    .S0(net465),
    .S1(net836),
    .X(net467));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(clknet_1_1__leaf_net178),
    .A1(clknet_1_1__leaf_net301),
    .A2(net803),
    .A3(net890),
    .S0(net907),
    .S1(net909),
    .X(net468));
 sky130_fd_sc_hd__mux4_1 c484 (.A0(net1182),
    .A1(net1100),
    .A2(net17),
    .A3(clknet_1_0__leaf_net289),
    .S0(net886),
    .S1(net904),
    .X(net469));
 sky130_fd_sc_hd__mux4_2 c485 (.A0(net977),
    .A1(clknet_1_0__leaf_net289),
    .A2(net378),
    .A3(net38),
    .S0(net1085),
    .S1(net1045),
    .X(net470));
 sky130_fd_sc_hd__mux4_1 c486 (.A0(net432),
    .A1(net390),
    .A2(net50),
    .A3(net345),
    .S0(net196),
    .S1(net1085),
    .X(net471));
 sky130_fd_sc_hd__mux4_1 c487 (.A0(net1019),
    .A1(net1010),
    .A2(net74),
    .A3(net390),
    .S0(clknet_1_1__leaf_net339),
    .S1(net812),
    .X(net472));
 sky130_fd_sc_hd__mux4_2 c488 (.A0(net17),
    .A1(net196),
    .A2(net1047),
    .A3(net1037),
    .S0(net890),
    .S1(net906),
    .X(net473));
 sky130_fd_sc_hd__mux4_1 c489 (.A0(net76),
    .A1(net1087),
    .A2(net54),
    .A3(net291),
    .S0(clknet_1_1__leaf_net339),
    .S1(net892),
    .X(net474));
 sky130_fd_sc_hd__xnor2_4 c49 (.A(net1107),
    .B(net39),
    .Y(net23));
 sky130_fd_sc_hd__mux4_1 c490 (.A0(net164),
    .A1(net1082),
    .A2(clknet_1_1__leaf_net174),
    .A3(clknet_1_1__leaf_net331),
    .S0(net183),
    .S1(net1092),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c491 (.A0(net197),
    .A1(net975),
    .A2(net1107),
    .A3(net404),
    .S0(net59),
    .S1(net910),
    .X(net476));
 sky130_fd_sc_hd__mux4_1 c492 (.A0(net292),
    .A1(net394),
    .A2(net59),
    .A3(net420),
    .S0(net1033),
    .S1(net404),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c493 (.A0(net344),
    .A1(net1002),
    .A2(net345),
    .A3(net166),
    .S0(net829),
    .S1(net910),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c494 (.A0(net468),
    .A1(net1009),
    .A2(net390),
    .A3(net378),
    .S0(clknet_1_1__leaf_net339),
    .S1(net905),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 c495 (.A0(net166),
    .A1(net1071),
    .A2(net1008),
    .A3(net394),
    .S0(net198),
    .S1(net1040),
    .X(net480));
 sky130_fd_sc_hd__mux4_1 c496 (.A0(net378),
    .A1(net166),
    .A2(net78),
    .A3(net393),
    .S0(net1079),
    .S1(clknet_1_0__leaf_net902),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 c497 (.A0(net452),
    .A1(clknet_1_0__leaf_net165),
    .A2(net477),
    .A3(net1034),
    .S0(net886),
    .S1(net911),
    .X(net482));
 sky130_fd_sc_hd__mux4_1 c498 (.A0(net475),
    .A1(net1045),
    .A2(net1165),
    .A3(net853),
    .S0(net906),
    .S1(net911),
    .X(net483));
 sky130_fd_sc_hd__mux4_1 c499 (.A0(clknet_1_0__leaf_net436),
    .A1(net481),
    .A2(net213),
    .A3(net1034),
    .S0(net1093),
    .S1(net905),
    .X(net484));
 sky130_fd_sc_hd__xnor2_4 c50 (.A(net1055),
    .B(net16),
    .Y(net24));
 sky130_fd_sc_hd__mux4_1 c500 (.A0(net74),
    .A1(net1035),
    .A2(net477),
    .A3(net1107),
    .S0(clknet_1_1__leaf_net177),
    .S1(net872),
    .X(net485));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(clknet_1_0__leaf_net456),
    .A1(net308),
    .A2(net285),
    .A3(net1034),
    .S0(net812),
    .S1(net848),
    .X(net486));
 sky130_fd_sc_hd__mux4_2 c502 (.A0(net308),
    .A1(net212),
    .A2(net38),
    .A3(net853),
    .S0(net872),
    .S1(net913),
    .X(net487));
 sky130_fd_sc_hd__mux4_1 c503 (.A0(net477),
    .A1(net139),
    .A2(clknet_1_0__leaf_net289),
    .A3(net465),
    .S0(net866),
    .S1(net913),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c504 (.A0(net441),
    .A1(clknet_1_0__leaf_net289),
    .A2(net125),
    .A3(net1036),
    .S0(net864),
    .S1(net913),
    .X(net489));
 sky130_fd_sc_hd__mux4_1 c505 (.A0(clknet_1_0__leaf_net289),
    .A1(clknet_1_0__leaf_net489),
    .A2(net60),
    .A3(clknet_1_1__leaf_net339),
    .S0(net910),
    .S1(net911),
    .X(net490));
 sky130_fd_sc_hd__mux4_1 c506 (.A0(net1019),
    .A1(net1050),
    .A2(net232),
    .A3(net159),
    .S0(net867),
    .S1(net914),
    .X(net491));
 sky130_fd_sc_hd__mux4_1 c507 (.A0(net60),
    .A1(clknet_1_1__leaf_net226),
    .A2(net1089),
    .A3(net285),
    .S0(net183),
    .S1(net866),
    .X(net492));
 sky130_fd_sc_hd__mux4_1 c508 (.A0(net1098),
    .A1(net354),
    .A2(net159),
    .A3(net1019),
    .S0(net1037),
    .S1(net1079),
    .X(net493));
 sky130_fd_sc_hd__mux4_1 c509 (.A0(clknet_1_0__leaf_net234),
    .A1(net1033),
    .A2(net1004),
    .A3(net76),
    .S0(net1008),
    .S1(net912),
    .X(net494));
 sky130_fd_sc_hd__xnor2_4 c51 (.A(net1083),
    .B(net1055),
    .Y(net25));
 sky130_fd_sc_hd__mux4_1 c510 (.A0(net355),
    .A1(net1039),
    .A2(net1019),
    .A3(net374),
    .S0(clknet_1_0__leaf_net470),
    .S1(net21),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 c511 (.A0(clknet_1_1__leaf_net352),
    .A1(net1138),
    .A2(net1004),
    .A3(net987),
    .S0(net1022),
    .S1(net207),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 c512 (.A0(net1009),
    .A1(net473),
    .A2(clknet_1_1__leaf_net496),
    .A3(clknet_1_0__leaf_net985),
    .S0(net795),
    .S1(net851),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 c513 (.A0(net492),
    .A1(clknet_1_0__leaf_net470),
    .A2(net13),
    .A3(net1021),
    .S0(net1009),
    .S1(net876),
    .X(net498));
 sky130_fd_sc_hd__mux4_1 c514 (.A0(net495),
    .A1(net210),
    .A2(net1034),
    .A3(net184),
    .S0(clknet_1_1__leaf_net222),
    .S1(net884),
    .X(net499));
 sky130_fd_sc_hd__mux4_2 c515 (.A0(net1025),
    .A1(net1019),
    .A2(clknet_1_1__leaf_net470),
    .A3(net1079),
    .S0(net851),
    .S1(net867),
    .X(net500));
 sky130_fd_sc_hd__mux4_1 c516 (.A0(net21),
    .A1(net229),
    .A2(net60),
    .A3(net473),
    .S0(net346),
    .S1(clknet_1_0__leaf_net496),
    .X(net501));
 sky130_fd_sc_hd__mux4_1 c517 (.A0(net159),
    .A1(clknet_1_0__leaf_net496),
    .A2(net1089),
    .A3(net876),
    .S0(net898),
    .S1(net915),
    .X(net502));
 sky130_fd_sc_hd__mux4_2 c518 (.A0(net210),
    .A1(net217),
    .A2(net207),
    .A3(net891),
    .S0(net916),
    .S1(net918),
    .X(net995));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net92),
    .A1(net100),
    .A2(net995),
    .A3(net1123),
    .S0(net895),
    .S1(net918),
    .X(net503));
 sky130_fd_sc_hd__a21bo_4 c52 (.A1(net16),
    .A2(net1095),
    .B1_N(net1047),
    .X(net26));
 sky130_fd_sc_hd__mux4_2 c520 (.A0(net346),
    .A1(net1036),
    .A2(net1030),
    .A3(clknet_1_0__leaf_net500),
    .S0(net795),
    .S1(net867),
    .X(net504));
 sky130_fd_sc_hd__mux4_1 c521 (.A0(clknet_1_1__leaf_net339),
    .A1(clknet_1_0__leaf_net504),
    .A2(net1099),
    .A3(clknet_1_1__leaf_net226),
    .S0(net873),
    .S1(net916),
    .X(net505));
 sky130_fd_sc_hd__mux4_1 c522 (.A0(net1030),
    .A1(clknet_1_1__leaf_net225),
    .A2(net995),
    .A3(clknet_1_1__leaf_net504),
    .S0(clknet_1_1__leaf_net234),
    .S1(net917),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 c523 (.A0(net1101),
    .A1(clknet_1_0__leaf_net504),
    .A2(net21),
    .A3(clknet_1_0__leaf_net499),
    .S0(net1022),
    .S1(net849),
    .X(net507));
 sky130_fd_sc_hd__mux4_1 c524 (.A0(net133),
    .A1(net473),
    .A2(net1105),
    .A3(net183),
    .S0(net808),
    .S1(net876),
    .X(net508));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(net374),
    .A1(net184),
    .A2(net285),
    .A3(net508),
    .S0(net866),
    .S1(net874),
    .X(net509));
 sky130_fd_sc_hd__mux4_1 c526 (.A0(net285),
    .A1(net508),
    .A2(net1087),
    .A3(net509),
    .S0(net978),
    .S1(net765),
    .X(net510));
 sky130_fd_sc_hd__mux4_2 c527 (.A0(clknet_1_1__leaf_net231),
    .A1(clknet_1_1__leaf_net351),
    .A2(net509),
    .A3(clknet_1_1__leaf_net504),
    .S0(net847),
    .S1(net915),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c528 (.A0(net386),
    .A1(net256),
    .A2(net391),
    .A3(net388),
    .S0(net385),
    .S1(net965),
    .X(net512));
 sky130_fd_sc_hd__xnor2_2 c529 (.A(net1090),
    .B(net396),
    .Y(net513));
 sky130_fd_sc_hd__a21bo_4 c53 (.A1(net22),
    .A2(net4),
    .B1_N(net1047),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 c530 (.A(net775),
    .X(net514));
 sky130_fd_sc_hd__a21bo_2 c531 (.A1(net1095),
    .A2(net240),
    .B1_N(net235),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_4 c532 (.A(net816),
    .X(net516));
 sky130_fd_sc_hd__xnor2_4 c533 (.A(net1088),
    .B(net516),
    .Y(net517));
 sky130_fd_sc_hd__dlymetal6s2s_1 c534 (.A(net816),
    .X(net989));
 sky130_fd_sc_hd__mux4_1 c535 (.A0(net514),
    .A1(net384),
    .A2(net1016),
    .A3(net257),
    .S0(net1066),
    .S1(net1068),
    .X(net518));
 sky130_fd_sc_hd__dlymetal6s2s_1 c536 (.A(net815),
    .X(net519));
 sky130_fd_sc_hd__a21bo_1 c537 (.A1(net380),
    .A2(net1070),
    .B1_N(net984),
    .X(net520));
 sky130_fd_sc_hd__xnor2_4 c538 (.A(net1118),
    .B(net517),
    .Y(net521));
 sky130_fd_sc_hd__a21bo_2 c539 (.A1(net968),
    .A2(net514),
    .B1_N(net235),
    .X(net522));
 sky130_fd_sc_hd__xnor2_4 c54 (.A(net11),
    .B(net1165),
    .Y(net28));
 sky130_fd_sc_hd__xnor2_2 c540 (.A(net522),
    .B(net1016),
    .Y(net523));
 sky130_fd_sc_hd__clkbuf_2 c541 (.A(net775),
    .X(net524));
 sky130_fd_sc_hd__xnor2_2 c542 (.A(net523),
    .B(net515),
    .Y(net525));
 sky130_fd_sc_hd__clkbuf_1 c543 (.A(net800),
    .X(net526));
 sky130_fd_sc_hd__a21bo_2 c544 (.A1(net235),
    .A2(net526),
    .B1_N(net517),
    .X(net527));
 sky130_fd_sc_hd__buf_1 c545 (.A(net815),
    .X(net528));
 sky130_fd_sc_hd__sdfbbn_1 c546 (.CLK_N(clknet_4_13_0_clk),
    .D(net524),
    .RESET_B(net527),
    .SCD(net528),
    .SCE(net1007),
    .SET_B(net382),
    .Q(net530),
    .Q_N(net529));
 sky130_fd_sc_hd__mux4_1 c547 (.A0(net523),
    .A1(net252),
    .A2(net527),
    .A3(net1007),
    .S0(net242),
    .S1(net919),
    .X(net531));
 sky130_fd_sc_hd__sdfbbn_1 c548 (.CLK_N(clknet_4_15_0_clk),
    .D(net1159),
    .RESET_B(net527),
    .SCD(net1007),
    .SCE(net516),
    .SET_B(net775),
    .Q(net533),
    .Q_N(net532));
 sky130_fd_sc_hd__sdfbbp_1 c549 (.CLK(clknet_4_15_0_clk),
    .D(net254),
    .RESET_B(net1066),
    .SCD(net528),
    .SCE(net533),
    .SET_B(net529),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__xnor2_4 c55 (.A(net27),
    .B(net17),
    .Y(net29));
 sky130_fd_sc_hd__a21bo_1 c550 (.A1(net1098),
    .A2(net398),
    .B1_N(net141),
    .X(net536));
 sky130_fd_sc_hd__a21bo_1 c551 (.A1(net262),
    .A2(net1163),
    .B1_N(net1078),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 c552 (.A(net770),
    .X(net1003));
 sky130_fd_sc_hd__a21bo_1 c553 (.A1(net383),
    .A2(net131),
    .B1_N(net812),
    .X(net538));
 sky130_fd_sc_hd__a31o_2 c554 (.A1(net383),
    .A2(net1086),
    .A3(net1040),
    .B1(net1064),
    .X(net539));
 sky130_fd_sc_hd__a21bo_1 c555 (.A1(net107),
    .A2(net524),
    .B1_N(net828),
    .X(net540));
 sky130_fd_sc_hd__sdfbbn_2 c556 (.CLK_N(clknet_4_13_0_clk),
    .D(net274),
    .RESET_B(net540),
    .SCD(net539),
    .SCE(net827),
    .SET_B(net919),
    .Q(net998),
    .Q_N(net541));
 sky130_fd_sc_hd__sdfrtp_1 c557 (.CLK(clknet_4_13_0_clk),
    .D(net526),
    .RESET_B(net1156),
    .SCD(net1064),
    .SCE(net400),
    .Q(net542));
 sky130_fd_sc_hd__clkbuf_1 c558 (.A(net770),
    .X(net543));
 sky130_fd_sc_hd__a41o_1 c559 (.A1(net528),
    .A2(net543),
    .A3(net406),
    .A4(net521),
    .B1(net1078),
    .X(net544));
 sky130_fd_sc_hd__a21bo_4 c56 (.A1(net25),
    .A2(net29),
    .B1_N(net26),
    .X(net30));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(net412),
    .A1(net544),
    .A2(net1157),
    .A3(net102),
    .S0(net1068),
    .S1(net1064),
    .X(net545));
 sky130_fd_sc_hd__buf_1 c561 (.A(net770),
    .X(net546));
 sky130_fd_sc_hd__buf_1 c562 (.A(net770),
    .X(net547));
 sky130_fd_sc_hd__mux4_1 c563 (.A0(net517),
    .A1(net401),
    .A2(net536),
    .A3(net539),
    .S0(net13),
    .S1(net1064),
    .X(net548));
 sky130_fd_sc_hd__buf_1 c564 (.A(net800),
    .X(net549));
 sky130_fd_sc_hd__mux4_1 c565 (.A0(net415),
    .A1(net546),
    .A2(net536),
    .A3(net403),
    .S0(net517),
    .S1(net1077),
    .X(net550));
 sky130_fd_sc_hd__mux4_2 c566 (.A0(net1157),
    .A1(net524),
    .A2(net519),
    .A3(net107),
    .S0(net404),
    .S1(net1070),
    .X(net551));
 sky130_fd_sc_hd__buf_1 c567 (.A(net797),
    .X(net552));
 sky130_fd_sc_hd__mux4_2 c568 (.A0(net519),
    .A1(net542),
    .A2(net539),
    .A3(net1064),
    .S0(net552),
    .S1(net920),
    .X(net997));
 sky130_fd_sc_hd__a41o_2 c569 (.A1(net546),
    .A2(net551),
    .A3(net552),
    .A4(net1064),
    .B1(net921),
    .X(net553));
 sky130_fd_sc_hd__xnor2_4 c57 (.A(net9),
    .B(net1051),
    .Y(net31));
 sky130_fd_sc_hd__a41o_2 c570 (.A1(net552),
    .A2(net997),
    .A3(net549),
    .A4(net553),
    .B1(net921),
    .X(net554));
 sky130_fd_sc_hd__mux4_2 c571 (.A0(net1084),
    .A1(net519),
    .A2(net997),
    .A3(net517),
    .S0(net554),
    .S1(net827),
    .X(net555));
 sky130_fd_sc_hd__mux4_2 c572 (.A0(net288),
    .A1(net530),
    .A2(net527),
    .A3(net975),
    .S0(net1064),
    .S1(net899),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 c573 (.A0(net131),
    .A1(clknet_1_1__leaf_net437),
    .A2(net1013),
    .A3(net828),
    .S0(clknet_1_0__leaf_net882),
    .S1(net921),
    .X(net557));
 sky130_fd_sc_hd__mux4_2 c574 (.A0(net384),
    .A1(net1110),
    .A2(net441),
    .A3(net1068),
    .S0(net828),
    .S1(net899),
    .X(net558));
 sky130_fd_sc_hd__mux4_1 c575 (.A0(net527),
    .A1(net1065),
    .A2(net555),
    .A3(net440),
    .S0(net1013),
    .S1(net1038),
    .X(net559));
 sky130_fd_sc_hd__mux4_1 c576 (.A0(net158),
    .A1(net1080),
    .A2(net255),
    .A3(net1088),
    .S0(net559),
    .S1(net920),
    .X(net560));
 sky130_fd_sc_hd__mux4_1 c577 (.A0(net407),
    .A1(net1042),
    .A2(net1014),
    .A3(net1013),
    .S0(net862),
    .S1(clknet_1_1__leaf_net901),
    .X(net561));
 sky130_fd_sc_hd__mux4_1 c578 (.A0(net133),
    .A1(net438),
    .A2(net989),
    .A3(net1038),
    .S0(net1076),
    .S1(clknet_1_1__leaf_net901),
    .X(net562));
 sky130_fd_sc_hd__mux4_1 c579 (.A0(net407),
    .A1(net133),
    .A2(net538),
    .A3(net287),
    .S0(net527),
    .S1(net1078),
    .X(net563));
 sky130_fd_sc_hd__xnor2_4 c58 (.A(net28),
    .B(net17),
    .Y(net32));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net1086),
    .A1(net288),
    .A2(net273),
    .A3(clknet_1_0__leaf_net561),
    .S0(net1013),
    .S1(net558),
    .X(net564));
 sky130_fd_sc_hd__mux4_1 c581 (.A0(net1110),
    .A1(net559),
    .A2(net240),
    .A3(clknet_1_0__leaf_net447),
    .S0(net1013),
    .S1(net921),
    .X(net565));
 sky130_fd_sc_hd__mux4_1 c582 (.A0(net563),
    .A1(clknet_1_0__leaf_net561),
    .A2(net1105),
    .A3(net553),
    .S0(clknet_1_1__leaf_net901),
    .S1(clknet_1_0__leaf_net922),
    .X(net566));
 sky130_fd_sc_hd__mux4_1 c583 (.A0(net549),
    .A1(net418),
    .A2(clknet_1_0__leaf_net562),
    .A3(net527),
    .S0(net30),
    .S1(net975),
    .X(net567));
 sky130_fd_sc_hd__mux4_1 c584 (.A0(net240),
    .A1(net25),
    .A2(net388),
    .A3(net404),
    .S0(net125),
    .S1(net1087),
    .X(net568));
 sky130_fd_sc_hd__mux4_1 c585 (.A0(net559),
    .A1(net149),
    .A2(clknet_1_0__leaf_net561),
    .A3(net287),
    .S0(net1013),
    .S1(net262),
    .X(net569));
 sky130_fd_sc_hd__mux4_1 c586 (.A0(net404),
    .A1(net515),
    .A2(net438),
    .A3(net1090),
    .S0(clknet_1_1__leaf_net567),
    .S1(clknet_1_0__leaf_net924),
    .X(net570));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_0__leaf_net570),
    .A1(net1013),
    .A2(net1095),
    .A3(net1009),
    .S0(net878),
    .S1(clknet_1_1__leaf_net924),
    .X(net571));
 sky130_fd_sc_hd__mux4_1 c588 (.A0(net515),
    .A1(net525),
    .A2(clknet_1_1__leaf_net570),
    .A3(net384),
    .S0(clknet_1_1__leaf_net301),
    .S1(clknet_1_1__leaf_net924),
    .X(net572));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net273),
    .A1(net398),
    .A2(net556),
    .A3(net1007),
    .S0(net554),
    .S1(clknet_1_1__leaf_net922),
    .X(net573));
 sky130_fd_sc_hd__a31o_1 c59 (.A1(net26),
    .A2(net9),
    .A3(net32),
    .B1(net1047),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 c590 (.A0(net384),
    .A1(net554),
    .A2(net407),
    .A3(clknet_1_0__leaf_net922),
    .S0(clknet_1_0__leaf_net924),
    .S1(net926),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c591 (.A0(net379),
    .A1(net427),
    .A2(net434),
    .A3(net1065),
    .S0(net817),
    .S1(net828),
    .X(net575));
 sky130_fd_sc_hd__mux4_1 c592 (.A0(net150),
    .A1(net558),
    .A2(net515),
    .A3(clknet_1_1__leaf_net574),
    .S0(net556),
    .S1(clknet_1_0__leaf_net924),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(clknet_1_0__leaf_net570),
    .A1(net556),
    .A2(net817),
    .A3(clknet_1_1__leaf_net881),
    .S0(net920),
    .S1(net925),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c594 (.A0(net400),
    .A1(net237),
    .A2(net1065),
    .A3(net1009),
    .S0(net1001),
    .S1(clknet_1_0__leaf_net903),
    .X(net578));
 sky130_fd_sc_hd__mux4_1 c595 (.A0(net13),
    .A1(net440),
    .A2(clknet_1_0__leaf_net315),
    .A3(net1093),
    .S0(net878),
    .S1(clknet_1_0__leaf_net903),
    .X(net579));
 sky130_fd_sc_hd__mux4_1 c596 (.A0(net259),
    .A1(net31),
    .A2(clknet_1_1__leaf_net174),
    .A3(net1096),
    .S0(clknet_1_1__leaf_net320),
    .S1(net1070),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c597 (.A0(net402),
    .A1(net1139),
    .A2(clknet_1_1__leaf_net313),
    .A3(net31),
    .S0(net1059),
    .S1(net1050),
    .X(net581));
 sky130_fd_sc_hd__mux4_1 c598 (.A0(net453),
    .A1(net1059),
    .A2(net1031),
    .A3(net1106),
    .S0(net841),
    .S1(net904),
    .X(net582));
 sky130_fd_sc_hd__mux4_2 c599 (.A0(net263),
    .A1(net127),
    .A2(net516),
    .A3(net148),
    .S0(net925),
    .S1(net930),
    .X(net583));
 sky130_fd_sc_hd__xnor2_4 c60 (.A(net1038),
    .B(net1047),
    .Y(net34));
 sky130_fd_sc_hd__mux4_1 c600 (.A0(net144),
    .A1(net1105),
    .A2(net184),
    .A3(net16),
    .S0(net888),
    .S1(net930),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 c601 (.A0(net1031),
    .A1(net1069),
    .A2(net583),
    .A3(net541),
    .S0(net402),
    .S1(net862),
    .X(net585));
 sky130_fd_sc_hd__mux4_1 c602 (.A0(net466),
    .A1(clknet_1_1__leaf_net178),
    .A2(clknet_1_1__leaf_net985),
    .A3(net127),
    .S0(net248),
    .S1(net930),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 c603 (.A0(net516),
    .A1(clknet_1_1__leaf_net301),
    .A2(clknet_1_1__leaf_net574),
    .A3(net1088),
    .S0(net1087),
    .S1(net931),
    .X(net587));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(net248),
    .A1(net1001),
    .A2(net1085),
    .A3(net860),
    .S0(net930),
    .S1(net932),
    .X(net588));
 sky130_fd_sc_hd__mux4_1 c605 (.A0(net247),
    .A1(clknet_1_0__leaf_net437),
    .A2(net588),
    .A3(net863),
    .S0(clknet_1_1__leaf_net881),
    .S1(net931),
    .X(net589));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net1093),
    .A1(net1098),
    .A2(net258),
    .A3(net931),
    .S0(net932),
    .S1(net933),
    .X(net590));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net16),
    .A1(net144),
    .A2(net583),
    .A3(net853),
    .S0(net932),
    .S1(net934),
    .X(net591));
 sky130_fd_sc_hd__mux4_1 c608 (.A0(net524),
    .A1(net525),
    .A2(clknet_1_1__leaf_net177),
    .A3(clknet_1_1__leaf_net178),
    .S0(net928),
    .S1(net934),
    .X(net592));
 sky130_fd_sc_hd__mux4_1 c609 (.A0(clknet_1_1__leaf_net315),
    .A1(net446),
    .A2(net843),
    .A3(clknet_1_0__leaf_net901),
    .S0(net933),
    .S1(net935),
    .X(net593));
 sky130_fd_sc_hd__a21bo_4 c61 (.A1(net32),
    .A2(net28),
    .B1_N(net1037),
    .X(net35));
 sky130_fd_sc_hd__mux4_1 c610 (.A0(net544),
    .A1(net157),
    .A2(net463),
    .A3(net466),
    .S0(net930),
    .S1(net934),
    .X(net594));
 sky130_fd_sc_hd__mux4_1 c611 (.A0(net1105),
    .A1(net184),
    .A2(clknet_1_1__leaf_net858),
    .A3(net928),
    .S0(net934),
    .S1(net935),
    .X(net595));
 sky130_fd_sc_hd__mux4_1 c612 (.A0(net1036),
    .A1(net38),
    .A2(net841),
    .A3(clknet_1_0__leaf_net901),
    .S0(net933),
    .S1(net934),
    .X(net596));
 sky130_fd_sc_hd__mux4_1 c613 (.A0(net30),
    .A1(clknet_1_0__leaf_net858),
    .A2(net931),
    .A3(net932),
    .S0(net933),
    .S1(net934),
    .X(net597));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net594),
    .A1(clknet_1_1__leaf_net597),
    .A2(net263),
    .A3(clknet_1_0__leaf_net596),
    .S0(clknet_1_0__leaf_net858),
    .S1(net934),
    .X(net598));
 sky130_fd_sc_hd__mux4_1 c615 (.A0(net1094),
    .A1(net30),
    .A2(net594),
    .A3(net588),
    .S0(net863),
    .S1(net937),
    .X(net599));
 sky130_fd_sc_hd__mux4_1 c616 (.A0(net588),
    .A1(net237),
    .A2(net134),
    .A3(net404),
    .S0(clknet_1_1__leaf_net177),
    .S1(net1125),
    .X(net600));
 sky130_fd_sc_hd__mux4_1 c617 (.A0(clknet_1_1__leaf_net489),
    .A1(net524),
    .A2(net525),
    .A3(net59),
    .S0(net487),
    .S1(net1117),
    .X(net601));
 sky130_fd_sc_hd__mux4_1 c618 (.A0(net1139),
    .A1(net487),
    .A2(clknet_1_1__leaf_net489),
    .A3(net1008),
    .S0(net399),
    .S1(net933),
    .X(net602));
 sky130_fd_sc_hd__mux4_1 c619 (.A0(net1107),
    .A1(net148),
    .A2(net1050),
    .A3(net446),
    .S0(net1061),
    .S1(net929),
    .X(net603));
 sky130_fd_sc_hd__a21bo_2 c62 (.A1(net1107),
    .A2(net35),
    .B1_N(net32),
    .X(net36));
 sky130_fd_sc_hd__mux4_1 c620 (.A0(net463),
    .A1(net1032),
    .A2(net1058),
    .A3(net975),
    .S0(clknet_1_0__leaf_net489),
    .S1(net237),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c621 (.A0(net38),
    .A1(clknet_1_0__leaf_net469),
    .A2(net1034),
    .A3(clknet_1_0__leaf_net489),
    .S0(net139),
    .S1(net905),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 c622 (.A0(clknet_1_0__leaf_net203),
    .A1(clknet_1_0__leaf_net313),
    .A2(net446),
    .A3(net404),
    .S0(net1059),
    .S1(net864),
    .X(net606));
 sky130_fd_sc_hd__mux4_1 c623 (.A0(net148),
    .A1(clknet_1_0__leaf_net595),
    .A2(net78),
    .A3(net907),
    .S0(net933),
    .S1(net938),
    .X(net607));
 sky130_fd_sc_hd__mux4_1 c624 (.A0(net136),
    .A1(clknet_1_0__leaf_net604),
    .A2(net1048),
    .A3(net848),
    .S0(net850),
    .S1(net872),
    .X(net608));
 sky130_fd_sc_hd__mux4_1 c625 (.A0(clknet_1_1__leaf_net469),
    .A1(net125),
    .A2(clknet_1_1__leaf_net489),
    .A3(net13),
    .S0(net963),
    .S1(net872),
    .X(net609));
 sky130_fd_sc_hd__mux4_1 c626 (.A0(clknet_1_0__leaf_net574),
    .A1(net538),
    .A2(clknet_1_1__leaf_net607),
    .A3(clknet_1_1__leaf_net203),
    .S0(net446),
    .S1(clknet_1_0__leaf_net881),
    .X(net610));
 sky130_fd_sc_hd__mux4_1 c627 (.A0(net1088),
    .A1(net1059),
    .A2(net441),
    .A3(clknet_1_0__leaf_net597),
    .S0(net1087),
    .S1(net845),
    .X(net611));
 sky130_fd_sc_hd__mux4_1 c628 (.A0(net25),
    .A1(clknet_1_0__leaf_net605),
    .A2(net608),
    .A3(net1013),
    .S0(clknet_1_0__leaf_net604),
    .S1(net487),
    .X(net612));
 sky130_fd_sc_hd__mux4_1 c629 (.A0(net441),
    .A1(net476),
    .A2(net1002),
    .A3(net434),
    .S0(clknet_1_1__leaf_net597),
    .S1(clknet_1_0__leaf_net469),
    .X(net613));
 sky130_fd_sc_hd__mux4_2 c63 (.A0(net36),
    .A1(net976),
    .A2(net23),
    .A3(net25),
    .S0(net1035),
    .S1(net975),
    .X(net37));
 sky130_fd_sc_hd__mux4_1 c630 (.A0(net1011),
    .A1(clknet_1_1__leaf_net174),
    .A2(clknet_1_1__leaf_net604),
    .A3(net125),
    .S0(net1050),
    .S1(clknet_1_1__leaf_net600),
    .X(net614));
 sky130_fd_sc_hd__mux4_1 c631 (.A0(net525),
    .A1(clknet_1_1__leaf_net177),
    .A2(net476),
    .A3(clknet_1_0__leaf_net881),
    .S0(net929),
    .S1(net933),
    .X(net615));
 sky130_fd_sc_hd__mux4_1 c632 (.A0(net404),
    .A1(clknet_1_0__leaf_net574),
    .A2(net998),
    .A3(clknet_1_0__leaf_net611),
    .S0(net237),
    .S1(net1000),
    .X(net616));
 sky130_fd_sc_hd__mux4_1 c633 (.A0(net1066),
    .A1(clknet_1_1__leaf_net605),
    .A2(clknet_1_1__leaf_net469),
    .A3(clknet_1_1__leaf_net822),
    .S0(net845),
    .S1(net850),
    .X(net617));
 sky130_fd_sc_hd__mux4_1 c634 (.A0(net617),
    .A1(clknet_1_1__leaf_net203),
    .A2(clknet_1_0__leaf_net609),
    .A3(net237),
    .S0(net865),
    .S1(net930),
    .X(net618));
 sky130_fd_sc_hd__a31o_1 c635 (.A1(net992),
    .A2(net850),
    .A3(net860),
    .B1(net869),
    .X(net619));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net239),
    .A1(net603),
    .A2(net59),
    .A3(net538),
    .S0(net832),
    .S1(net868),
    .X(net620));
 sky130_fd_sc_hd__mux4_1 c637 (.A0(net620),
    .A1(net619),
    .A2(clknet_1_1__leaf_net609),
    .A3(clknet_1_0__leaf_net437),
    .S0(net855),
    .S1(clknet_1_1__leaf_net994),
    .X(net621));
 sky130_fd_sc_hd__mux4_2 c64 (.A0(net35),
    .A1(net30),
    .A2(net37),
    .A3(net1037),
    .S0(net1035),
    .S1(net1047),
    .X(net38));
 sky130_fd_sc_hd__mux4_1 c643 (.A0(clknet_1_1__leaf_net165),
    .A1(clknet_1_0__leaf_net313),
    .A2(net1066),
    .A3(net999),
    .S0(net847),
    .S1(net926),
    .X(net622));
 sky130_fd_sc_hd__mux4_1 c644 (.A0(net1073),
    .A1(net66),
    .A2(clknet_1_0__leaf_net221),
    .A3(net1103),
    .S0(net1041),
    .S1(net184),
    .X(net623));
 sky130_fd_sc_hd__mux4_1 c645 (.A0(net623),
    .A1(net139),
    .A2(clknet_1_0__leaf_net600),
    .A3(clknet_1_1__leaf_net165),
    .S0(net1094),
    .S1(clknet_1_1__leaf_net500),
    .X(net624));
 sky130_fd_sc_hd__mux4_1 c646 (.A0(net434),
    .A1(net1022),
    .A2(net558),
    .A3(net1033),
    .S0(clknet_1_1__leaf_net221),
    .S1(clknet_1_0__leaf_net994),
    .X(net625));
 sky130_fd_sc_hd__mux4_1 c647 (.A0(net1021),
    .A1(clknet_1_0__leaf_net320),
    .A2(clknet_1_0__leaf_net600),
    .A3(net834),
    .S0(net864),
    .S1(net866),
    .X(net626));
 sky130_fd_sc_hd__a41o_1 c648 (.A1(net1008),
    .A2(net184),
    .A3(clknet_1_1__leaf_net165),
    .A4(net1006),
    .B1(clknet_1_0__leaf_net881),
    .X(net627));
 sky130_fd_sc_hd__mux4_1 c649 (.A0(net198),
    .A1(clknet_1_0__leaf_net313),
    .A2(net992),
    .A3(net995),
    .S0(net914),
    .S1(net939),
    .X(net628));
 sky130_fd_sc_hd__xnor2_4 c65 (.A(net1099),
    .B(net9),
    .Y(net39));
 sky130_fd_sc_hd__mux4_1 c650 (.A0(clknet_1_0__leaf_net607),
    .A1(net130),
    .A2(net1088),
    .A3(net864),
    .S0(net912),
    .S1(net918),
    .X(net1005));
 sky130_fd_sc_hd__mux4_1 c651 (.A0(clknet_1_0__leaf_net500),
    .A1(net1105),
    .A2(net137),
    .A3(net1073),
    .S0(net817),
    .S1(net914),
    .X(net629));
 sky130_fd_sc_hd__mux4_1 c652 (.A0(net1037),
    .A1(net232),
    .A2(net622),
    .A3(net1021),
    .S0(net198),
    .S1(net912),
    .X(net630));
 sky130_fd_sc_hd__mux4_1 c653 (.A0(clknet_1_1__leaf_net499),
    .A1(clknet_1_0__leaf_net437),
    .A2(net1048),
    .A3(net1022),
    .S0(net100),
    .S1(net844),
    .X(net631));
 sky130_fd_sc_hd__mux4_1 c654 (.A0(net50),
    .A1(net100),
    .A2(clknet_1_1__leaf_net222),
    .A3(net1008),
    .S0(clknet_1_0__leaf_net881),
    .S1(net939),
    .X(net632));
 sky130_fd_sc_hd__mux4_1 c655 (.A0(net141),
    .A1(net995),
    .A2(clknet_1_0__leaf_net822),
    .A3(net841),
    .S0(net856),
    .S1(net891),
    .X(net633));
 sky130_fd_sc_hd__mux4_1 c656 (.A0(net633),
    .A1(net844),
    .A2(clknet_1_0__leaf_net881),
    .A3(net891),
    .S0(net917),
    .S1(net939),
    .X(net634));
 sky130_fd_sc_hd__mux4_1 c657 (.A0(net1089),
    .A1(clknet_1_0__leaf_net331),
    .A2(net510),
    .A3(net1043),
    .S0(net856),
    .S1(net939),
    .X(net635));
 sky130_fd_sc_hd__mux4_1 c658 (.A0(clknet_1_0__leaf_net635),
    .A1(net59),
    .A2(net1090),
    .A3(net841),
    .S0(net870),
    .S1(net939),
    .X(net996));
 sky130_fd_sc_hd__mux4_1 c659 (.A0(net629),
    .A1(clknet_1_0__leaf_net320),
    .A2(net628),
    .A3(clknet_1_1__leaf_net996),
    .S0(clknet_1_1__leaf_net635),
    .S1(net831),
    .X(net636));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net13),
    .B(net26),
    .Y(net1001));
 sky130_fd_sc_hd__a41o_2 c660 (.A1(net1106),
    .A2(net249),
    .A3(net963),
    .A4(net1107),
    .B1(net521),
    .X(net637));
 sky130_fd_sc_hd__xnor2_2 c661 (.A(net984),
    .B(net637),
    .Y(net638));
 sky130_fd_sc_hd__xnor2_2 c662 (.A(net396),
    .B(net1107),
    .Y(net639));
 sky130_fd_sc_hd__xnor2_1 c663 (.A(net1103),
    .B(net639),
    .Y(net640));
 sky130_fd_sc_hd__buf_1 c664 (.A(net768),
    .X(net641));
 sky130_fd_sc_hd__xnor2_1 c665 (.A(net1119),
    .B(net638),
    .Y(net642));
 sky130_fd_sc_hd__xnor2_2 c666 (.A(net513),
    .B(net641),
    .Y(net643));
 sky130_fd_sc_hd__buf_1 c667 (.A(net768),
    .X(net644));
 sky130_fd_sc_hd__xnor2_2 c668 (.A(net247),
    .B(net775),
    .Y(net645));
 sky130_fd_sc_hd__sdfbbn_1 c669 (.CLK_N(clknet_4_15_0_clk),
    .D(net1095),
    .RESET_B(net1007),
    .SCD(net645),
    .SCE(net1110),
    .SET_B(net1043),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__xnor2_4 c67 (.A(net1053),
    .B(net17),
    .Y(net40));
 sky130_fd_sc_hd__xnor2_2 c670 (.A(net647),
    .B(net522),
    .Y(net648));
 sky130_fd_sc_hd__xnor2_2 c671 (.A(net648),
    .B(net643),
    .Y(net649));
 sky130_fd_sc_hd__xnor2_1 c672 (.A(net639),
    .B(net971),
    .Y(net650));
 sky130_fd_sc_hd__dlymetal6s2s_1 c673 (.A(net797),
    .X(net651));
 sky130_fd_sc_hd__a21bo_1 c674 (.A1(net641),
    .A2(net385),
    .B1_N(net648),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_2 c675 (.A(net1162),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 c676 (.A(net768),
    .X(net654));
 sky130_fd_sc_hd__a21bo_1 c677 (.A1(net521),
    .A2(net1119),
    .B1_N(net1069),
    .X(net655));
 sky130_fd_sc_hd__a41o_2 c678 (.A1(net651),
    .A2(net655),
    .A3(net247),
    .A4(net249),
    .B1(net522),
    .X(net656));
 sky130_fd_sc_hd__a41o_2 c679 (.A1(net522),
    .A2(net648),
    .A3(net641),
    .A4(net654),
    .B1(net970),
    .X(net657));
 sky130_fd_sc_hd__xnor2_4 c68 (.A(net18),
    .B(net1046),
    .Y(net41));
 sky130_fd_sc_hd__mux4_1 c680 (.A0(net654),
    .A1(net249),
    .A2(net655),
    .A3(net639),
    .S0(net657),
    .S1(net645),
    .X(net658));
 sky130_fd_sc_hd__sdfbbp_1 c681 (.CLK(clknet_4_15_0_clk),
    .D(net645),
    .RESET_B(net657),
    .SCD(net520),
    .SCE(net989),
    .SET_B(net1151),
    .Q(net660),
    .Q_N(net659));
 sky130_fd_sc_hd__a41o_1 c682 (.A1(net533),
    .A2(net653),
    .A3(net1009),
    .A4(net1069),
    .B1(net1155),
    .X(net661));
 sky130_fd_sc_hd__sdfbbn_2 c683 (.CLK_N(clknet_4_15_0_clk),
    .D(net639),
    .RESET_B(net638),
    .SCD(net637),
    .SCE(net405),
    .SET_B(net657),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__mux4_1 c684 (.A0(net655),
    .A1(net647),
    .A2(net657),
    .A3(net1069),
    .S0(net417),
    .S1(net551),
    .X(net664));
 sky130_fd_sc_hd__a31o_1 c685 (.A1(net535),
    .A2(net645),
    .A3(net1103),
    .B1(net1076),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 c686 (.A0(net539),
    .A1(net640),
    .A2(net1071),
    .A3(net1069),
    .S0(net534),
    .S1(net1076),
    .X(net666));
 sky130_fd_sc_hd__a41o_1 c687 (.A1(net656),
    .A2(net417),
    .A3(net967),
    .A4(net1069),
    .B1(net761),
    .X(net667));
 sky130_fd_sc_hd__a31o_1 c688 (.A1(net533),
    .A2(net663),
    .A3(net539),
    .B1(net831),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 c689 (.A0(net547),
    .A1(net663),
    .A2(net657),
    .A3(net1010),
    .S0(net1098),
    .S1(net827),
    .X(net669));
 sky130_fd_sc_hd__xnor2_2 c69 (.A(net972),
    .B(net1072),
    .Y(net42));
 sky130_fd_sc_hd__a41o_1 c690 (.A1(net645),
    .A2(net659),
    .A3(net662),
    .A4(net646),
    .B1(net760),
    .X(net670));
 sky130_fd_sc_hd__a31o_1 c691 (.A1(net406),
    .A2(net535),
    .A3(net1064),
    .B1(net385),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net640),
    .A1(net1126),
    .A2(net1107),
    .A3(net662),
    .S0(net1053),
    .S1(net1010),
    .X(net672));
 sky130_fd_sc_hd__a41o_1 c693 (.A1(net638),
    .A2(net1093),
    .A3(net532),
    .A4(net2),
    .B1(net108),
    .X(net673));
 sky130_fd_sc_hd__a41o_1 c694 (.A1(net540),
    .A2(net420),
    .A3(net980),
    .A4(net537),
    .B1(net1158),
    .X(net674));
 sky130_fd_sc_hd__a41o_1 c695 (.A1(net419),
    .A2(net534),
    .A3(net662),
    .A4(net1165),
    .B1(net940),
    .X(net675));
 sky130_fd_sc_hd__mux4_1 c696 (.A0(net670),
    .A1(net663),
    .A2(net1080),
    .A3(net551),
    .S0(net812),
    .S1(net1077),
    .X(net676));
 sky130_fd_sc_hd__a41o_1 c697 (.A1(net673),
    .A2(net660),
    .A3(net521),
    .A4(net553),
    .B1(net1077),
    .X(net677));
 sky130_fd_sc_hd__a31o_1 c698 (.A1(net387),
    .A2(net141),
    .A3(net1069),
    .B1(net838),
    .X(net678));
 sky130_fd_sc_hd__a31o_1 c699 (.A1(net108),
    .A2(net1065),
    .A3(net761),
    .B1(net1077),
    .X(net679));
 sky130_fd_sc_hd__xnor2_4 c70 (.A(net1073),
    .B(net41),
    .Y(net988));
 sky130_fd_sc_hd__mux4_1 c700 (.A0(net679),
    .A1(net980),
    .A2(net662),
    .A3(net408),
    .S0(net1071),
    .S1(net865),
    .X(net680));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net387),
    .A1(net651),
    .A2(net532),
    .A3(net662),
    .S0(net1065),
    .S1(net1139),
    .X(net681));
 sky130_fd_sc_hd__a41o_1 c702 (.A1(net978),
    .A2(net539),
    .A3(net547),
    .A4(net796),
    .B1(net831),
    .X(net682));
 sky130_fd_sc_hd__a21bo_1 c703 (.A1(net682),
    .A2(net257),
    .B1_N(net679),
    .X(net683));
 sky130_fd_sc_hd__mux4_1 c704 (.A0(net1040),
    .A1(net1007),
    .A2(net663),
    .A3(net1139),
    .S0(net832),
    .S1(net1151),
    .X(net684));
 sky130_fd_sc_hd__mux4_1 c705 (.A0(net555),
    .A1(net401),
    .A2(net676),
    .A3(net659),
    .S0(net247),
    .S1(clknet_1_1__leaf_net882),
    .X(net685));
 sky130_fd_sc_hd__mux4_1 c706 (.A0(net683),
    .A1(net0),
    .A2(net1012),
    .A3(net521),
    .S0(net656),
    .S1(net970),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 c707 (.A0(net1007),
    .A1(net675),
    .A2(net127),
    .A3(net555),
    .S0(net1040),
    .S1(net941),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 c708 (.A0(net551),
    .A1(net405),
    .A2(net141),
    .A3(net649),
    .S0(net973),
    .S1(clknet_1_1__leaf_net923),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 c709 (.A0(net418),
    .A1(net670),
    .A2(clknet_1_1__leaf_net561),
    .A3(net1007),
    .S0(net800),
    .S1(clknet_1_1__leaf_net882),
    .X(net689));
 sky130_fd_sc_hd__xnor2_4 c71 (.A(net964),
    .B(net1146),
    .Y(net43));
 sky130_fd_sc_hd__mux4_2 c710 (.A0(net408),
    .A1(net1011),
    .A2(net657),
    .A3(net1007),
    .S0(net663),
    .S1(net1065),
    .X(net690));
 sky130_fd_sc_hd__mux4_1 c711 (.A0(net537),
    .A1(net1053),
    .A2(net1014),
    .A3(net257),
    .S0(net982),
    .S1(clknet_1_0__leaf_net942),
    .X(net691));
 sky130_fd_sc_hd__mux4_1 c712 (.A0(net530),
    .A1(net1110),
    .A2(net162),
    .A3(net1043),
    .S0(net1009),
    .S1(net657),
    .X(net692));
 sky130_fd_sc_hd__mux4_1 c713 (.A0(clknet_1_1__leaf_net567),
    .A1(net521),
    .A2(net1070),
    .A3(net656),
    .S0(net662),
    .S1(net899),
    .X(net693));
 sky130_fd_sc_hd__mux4_1 c714 (.A0(net660),
    .A1(net521),
    .A2(net3),
    .A3(net529),
    .S0(clknet_1_1__leaf_net567),
    .S1(net1069),
    .X(net694));
 sky130_fd_sc_hd__mux4_1 c715 (.A0(net405),
    .A1(clknet_1_1__leaf_net693),
    .A2(net521),
    .A3(net840),
    .S0(net865),
    .S1(clknet_1_1__leaf_net882),
    .X(net695));
 sky130_fd_sc_hd__mux4_1 c716 (.A0(net418),
    .A1(net965),
    .A2(net662),
    .A3(net796),
    .S0(net846),
    .S1(clknet_1_1__leaf_net944),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c717 (.A0(net537),
    .A1(net247),
    .A2(clknet_1_1__leaf_net694),
    .A3(net657),
    .S0(net828),
    .S1(clknet_1_1__leaf_net942),
    .X(net697));
 sky130_fd_sc_hd__mux4_1 c718 (.A0(net651),
    .A1(net420),
    .A2(net553),
    .A3(net427),
    .S0(net663),
    .S1(clknet_1_1__leaf_net944),
    .X(net698));
 sky130_fd_sc_hd__mux4_1 c719 (.A0(clknet_1_0__leaf_net447),
    .A1(net671),
    .A2(net427),
    .A3(net555),
    .S0(clknet_1_1__leaf_net694),
    .S1(net662),
    .X(net699));
 sky130_fd_sc_hd__xnor2_2 c72 (.A(net1106),
    .B(net18),
    .Y(net44));
 sky130_fd_sc_hd__mux4_1 c720 (.A0(clknet_1_1__leaf_net447),
    .A1(net158),
    .A2(net1058),
    .A3(net800),
    .S0(clknet_1_1__leaf_net882),
    .S1(net941),
    .X(net700));
 sky130_fd_sc_hd__mux4_1 c721 (.A0(clknet_1_1__leaf_net562),
    .A1(net649),
    .A2(clknet_1_1__leaf_net700),
    .A3(net683),
    .S0(net663),
    .S1(net941),
    .X(net701));
 sky130_fd_sc_hd__mux4_1 c722 (.A0(net158),
    .A1(clknet_1_0__leaf_net693),
    .A2(net649),
    .A3(net846),
    .S0(net945),
    .S1(net947),
    .X(net702));
 sky130_fd_sc_hd__mux4_1 c723 (.A0(net668),
    .A1(net554),
    .A2(net840),
    .A3(net843),
    .S0(clknet_1_1__leaf_net943),
    .S1(net947),
    .X(net703));
 sky130_fd_sc_hd__mux4_1 c724 (.A0(net657),
    .A1(net671),
    .A2(net840),
    .A3(net899),
    .S0(net946),
    .S1(net948),
    .X(net704));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net649),
    .A1(clknet_1_1__leaf_net561),
    .A2(net675),
    .A3(clknet_1_1__leaf_net703),
    .S0(net852),
    .S1(net949),
    .X(net705));
 sky130_fd_sc_hd__mux4_1 c726 (.A0(net1099),
    .A1(net1058),
    .A2(net554),
    .A3(net553),
    .S0(clknet_1_0__leaf_net596),
    .S1(net583),
    .X(net706));
 sky130_fd_sc_hd__mux4_1 c727 (.A0(net257),
    .A1(net583),
    .A2(net650),
    .A3(clknet_1_1__leaf_net315),
    .S0(net888),
    .S1(net927),
    .X(net707));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(net553),
    .A1(net668),
    .A2(net1014),
    .A3(net653),
    .S0(net948),
    .S1(net951),
    .X(net708));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(net960),
    .A1(clknet_1_0__leaf_net696),
    .A2(net283),
    .A3(net888),
    .S0(clknet_1_0__leaf_net942),
    .S1(net951),
    .X(net709));
 sky130_fd_sc_hd__a21bo_2 c73 (.A1(net23),
    .A2(net1089),
    .B1_N(net1),
    .X(net45));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net1065),
    .A1(net553),
    .A2(net852),
    .A3(net887),
    .S0(clknet_1_1__leaf_net903),
    .S1(clknet_1_0__leaf_net944),
    .X(net710));
 sky130_fd_sc_hd__mux4_1 c731 (.A0(net162),
    .A1(net666),
    .A2(net395),
    .A3(net971),
    .S0(clknet_1_0__leaf_net923),
    .S1(net950),
    .X(net711));
 sky130_fd_sc_hd__mux4_1 c732 (.A0(net149),
    .A1(net708),
    .A2(net650),
    .A3(net1095),
    .S0(net1035),
    .S1(net1077),
    .X(net712));
 sky130_fd_sc_hd__mux4_1 c733 (.A0(net650),
    .A1(net13),
    .A2(net710),
    .A3(net663),
    .S0(net257),
    .S1(net930),
    .X(net713));
 sky130_fd_sc_hd__mux4_1 c734 (.A0(clknet_1_1__leaf_net315),
    .A1(net1061),
    .A2(net1011),
    .A3(clknet_1_1__leaf_net596),
    .S0(net1058),
    .S1(net1066),
    .X(net714));
 sky130_fd_sc_hd__mux4_1 c735 (.A0(net680),
    .A1(net127),
    .A2(net1069),
    .A3(net1035),
    .S0(net991),
    .S1(net952),
    .X(net715));
 sky130_fd_sc_hd__mux4_1 c736 (.A0(net1149),
    .A1(net676),
    .A2(clknet_1_0__leaf_net700),
    .A3(net1053),
    .S0(clknet_1_1__leaf_net161),
    .S1(clknet_1_1__leaf_net942),
    .X(net716));
 sky130_fd_sc_hd__mux4_1 c737 (.A0(net2),
    .A1(net258),
    .A2(net1009),
    .A3(net1124),
    .S0(clknet_1_0__leaf_net709),
    .S1(net257),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c738 (.A0(net283),
    .A1(net963),
    .A2(clknet_1_1__leaf_net706),
    .A3(clknet_1_0__leaf_net923),
    .S0(net952),
    .S1(net953),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 c739 (.A0(net247),
    .A1(net1069),
    .A2(net665),
    .A3(net1071),
    .S0(clknet_1_1__leaf_net902),
    .S1(net952),
    .X(net719));
 sky130_fd_sc_hd__xnor2_4 c74 (.A(net976),
    .B(net1056),
    .Y(net46));
 sky130_fd_sc_hd__mux4_1 c740 (.A0(net458),
    .A1(net667),
    .A2(net978),
    .A3(net837),
    .S0(net849),
    .S1(net861),
    .X(net720));
 sky130_fd_sc_hd__mux4_1 c741 (.A0(clknet_1_0__leaf_net703),
    .A1(net149),
    .A2(net162),
    .A3(net837),
    .S0(clknet_1_0__leaf_net942),
    .S1(net952),
    .X(net721));
 sky130_fd_sc_hd__mux4_1 c742 (.A0(clknet_1_1__leaf_net596),
    .A1(net553),
    .A2(clknet_1_1__leaf_net721),
    .A3(net427),
    .S0(net986),
    .S1(net953),
    .X(net722));
 sky130_fd_sc_hd__mux4_1 c743 (.A0(net715),
    .A1(clknet_1_1__leaf_net696),
    .A2(net680),
    .A3(net668),
    .S0(net136),
    .S1(net952),
    .X(net723));
 sky130_fd_sc_hd__mux4_1 c744 (.A0(net666),
    .A1(net713),
    .A2(net644),
    .A3(net162),
    .S0(net948),
    .S1(net953),
    .X(net724));
 sky130_fd_sc_hd__mux4_1 c745 (.A0(net568),
    .A1(net723),
    .A2(net283),
    .A3(net399),
    .S0(net861),
    .S1(net954),
    .X(net725));
 sky130_fd_sc_hd__a41o_1 c746 (.A1(net1014),
    .A2(net832),
    .A3(clknet_1_0__leaf_net943),
    .A4(net954),
    .B1(net955),
    .X(net726));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(clknet_1_1__leaf_net709),
    .A1(net667),
    .A2(net726),
    .A3(net1065),
    .S0(net952),
    .S1(net955),
    .X(net727));
 sky130_fd_sc_hd__mux4_1 c748 (.A0(net644),
    .A1(net1165),
    .A2(net965),
    .A3(net1066),
    .S0(net637),
    .S1(net855),
    .X(net728));
 sky130_fd_sc_hd__mux4_1 c749 (.A0(clknet_1_0__leaf_net706),
    .A1(net637),
    .A2(net718),
    .A3(net1009),
    .S0(net1058),
    .S1(net1066),
    .X(net729));
 sky130_fd_sc_hd__xnor2_2 c75 (.A(net41),
    .B(net46),
    .Y(net47));
 sky130_fd_sc_hd__mux4_1 c750 (.A0(net1125),
    .A1(net136),
    .A2(clknet_1_1__leaf_net161),
    .A3(net831),
    .S0(net849),
    .S1(net957),
    .X(net730));
 sky130_fd_sc_hd__mux4_1 c751 (.A0(net213),
    .A1(net730),
    .A2(net78),
    .A3(clknet_1_1__leaf_net902),
    .S0(net951),
    .S1(net956),
    .X(net731));
 sky130_fd_sc_hd__mux4_1 c752 (.A0(net399),
    .A1(net427),
    .A2(net1124),
    .A3(net1012),
    .S0(clknet_1_1__leaf_net161),
    .S1(net952),
    .X(net732));
 sky130_fd_sc_hd__mux4_1 c753 (.A0(net975),
    .A1(net1071),
    .A2(net153),
    .A3(net987),
    .S0(net1035),
    .S1(clknet_1_0__leaf_net944),
    .X(net733));
 sky130_fd_sc_hd__mux4_1 c754 (.A0(net982),
    .A1(net1011),
    .A2(net1043),
    .A3(net803),
    .S0(net1164),
    .S1(net1154),
    .X(net734));
 sky130_fd_sc_hd__mux4_1 c755 (.A0(net731),
    .A1(net663),
    .A2(net1001),
    .A3(net136),
    .S0(net1058),
    .S1(net955),
    .X(net735));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(clknet_1_0__leaf_net609),
    .A1(net1011),
    .A2(clknet_1_0__leaf_net567),
    .A3(net786),
    .S0(net930),
    .S1(net938),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 c757 (.A0(net1059),
    .A1(clknet_1_0__leaf_net567),
    .A2(net982),
    .A3(net978),
    .S0(clknet_1_0__leaf_net694),
    .S1(net930),
    .X(net737));
 sky130_fd_sc_hd__mux4_1 c758 (.A0(clknet_1_0__leaf_net595),
    .A1(net54),
    .A2(net965),
    .A3(clknet_1_0__leaf_net721),
    .S0(net1099),
    .S1(net870),
    .X(net738));
 sky130_fd_sc_hd__mux4_1 c759 (.A0(clknet_1_0__leaf_net597),
    .A1(net465),
    .A2(net1165),
    .A3(net644),
    .S0(clknet_1_0__leaf_net611),
    .S1(net786),
    .X(net739));
 sky130_fd_sc_hd__xnor2_4 c76 (.A(net979),
    .B(net35),
    .Y(net48));
 sky130_fd_sc_hd__mux4_1 c760 (.A0(net34),
    .A1(net656),
    .A2(net78),
    .A3(net728),
    .S0(net987),
    .S1(net1012),
    .X(net740));
 sky130_fd_sc_hd__mux4_1 c761 (.A0(net554),
    .A1(clknet_1_0__leaf_net694),
    .A2(net719),
    .A3(net1011),
    .S0(net1066),
    .S1(net952),
    .X(net741));
 sky130_fd_sc_hd__mux4_1 c762 (.A0(net733),
    .A1(net665),
    .A2(net554),
    .A3(net907),
    .S0(net957),
    .S1(net958),
    .X(net742));
 sky130_fd_sc_hd__mux4_1 c763 (.A0(net1013),
    .A1(clknet_1_0__leaf_net721),
    .A2(net738),
    .A3(net1066),
    .S0(net872),
    .S1(net936),
    .X(net743));
 sky130_fd_sc_hd__mux4_1 c764 (.A0(net1093),
    .A1(net1087),
    .A2(net739),
    .A3(net1013),
    .S0(net852),
    .S1(net871),
    .X(net744));
 sky130_fd_sc_hd__mux4_1 c765 (.A0(net134),
    .A1(net1012),
    .A2(net420),
    .A3(net742),
    .S0(net137),
    .S1(clknet_1_1__leaf_net595),
    .X(net745));
 sky130_fd_sc_hd__mux4_1 c766 (.A0(net153),
    .A1(net969),
    .A2(net743),
    .A3(net246),
    .S0(net840),
    .S1(clknet_1_1__leaf_net994),
    .X(net746));
 sky130_fd_sc_hd__mux4_1 c767 (.A0(clknet_1_1__leaf_net161),
    .A1(net744),
    .A2(net1048),
    .A3(clknet_1_1__leaf_net858),
    .S0(net869),
    .S1(net936),
    .X(net747));
 sky130_fd_sc_hd__mux4_1 c768 (.A0(net653),
    .A1(net137),
    .A2(clknet_1_1__leaf_net611),
    .A3(net865),
    .S0(net871),
    .S1(net907),
    .X(net748));
 sky130_fd_sc_hd__mux4_1 c769 (.A0(net965),
    .A1(net748),
    .A2(net849),
    .A3(net853),
    .S0(net956),
    .S1(net959));
 sky130_fd_sc_hd__xnor2_2 c77 (.A(net46),
    .B(net964),
    .Y(net993));
 sky130_fd_sc_hd__xnor2_2 c78 (.A(net1101),
    .B(net1056),
    .Y(net49));
 sky130_fd_sc_hd__a21bo_2 c79 (.A1(net1046),
    .A2(net45),
    .B1_N(net49),
    .X(net50));
 sky130_fd_sc_hd__a41o_2 c80 (.A1(net976),
    .A2(net47),
    .A3(net49),
    .A4(net1073),
    .B1(net26),
    .X(net51));
 sky130_fd_sc_hd__xnor2_2 c81 (.A(net18),
    .B(net1083),
    .Y(net52));
 sky130_fd_sc_hd__a41o_2 c82 (.A1(net12),
    .A2(net1055),
    .A3(net1041),
    .A4(net1046),
    .B1(net39),
    .X(net53));
 sky130_fd_sc_hd__xnor2_4 c83 (.A(net1041),
    .B(net53),
    .Y(net54));
 sky130_fd_sc_hd__mux4_2 c84 (.A0(net43),
    .A1(net1041),
    .A2(net54),
    .A3(net48),
    .S0(net45),
    .S1(net51),
    .X(net55));
 sky130_fd_sc_hd__xnor2_2 c85 (.A(net49),
    .B(net43),
    .Y(net56));
 sky130_fd_sc_hd__mux4_2 c86 (.A0(net54),
    .A1(net56),
    .A2(net1031),
    .A3(net1046),
    .S0(net18),
    .S1(net979),
    .X(net57));
 sky130_fd_sc_hd__mux4_2 c87 (.A0(net47),
    .A1(net56),
    .A2(net36),
    .A3(net988),
    .S0(net57),
    .S1(net1031),
    .X(net58));
 sky130_fd_sc_hd__a31o_4 c88 (.A1(net1035),
    .A2(net1060),
    .A3(net12),
    .B1(net32),
    .X(net59));
 sky130_fd_sc_hd__xnor2_4 c89 (.A(net1049),
    .B(net59),
    .Y(net60));
 sky130_fd_sc_hd__xnor2_4 c90 (.A(net11),
    .B(net35),
    .Y(net987));
 sky130_fd_sc_hd__xnor2_2 c91 (.A(net35),
    .B(net1048),
    .Y(net61));
 sky130_fd_sc_hd__xnor2_4 c92 (.A(net1062),
    .B(net1085),
    .Y(net62));
 sky130_fd_sc_hd__a21bo_1 c93 (.A1(net25),
    .A2(net32),
    .B1_N(net1073),
    .X(net63));
 sky130_fd_sc_hd__a41o_1 c94 (.A1(net1092),
    .A2(net61),
    .A3(net62),
    .A4(net63),
    .B1(net60),
    .X(net64));
 sky130_fd_sc_hd__xnor2_2 c95 (.A(net47),
    .B(net62),
    .Y(net65));
 sky130_fd_sc_hd__a31o_1 c96 (.A1(net1061),
    .A2(net18),
    .A3(net65),
    .B1(net53),
    .X(net66));
 sky130_fd_sc_hd__a21bo_2 c97 (.A1(net1091),
    .A2(net61),
    .B1_N(net1047),
    .X(net67));
 sky130_fd_sc_hd__a21bo_1 c98 (.A1(net63),
    .A2(net54),
    .B1_N(net41),
    .X(net68));
 sky130_fd_sc_hd__a31o_1 c99 (.A1(net65),
    .A2(net67),
    .A3(net988),
    .B1(net60),
    .X(net69));
 sky130_fd_sc_hd__a31o_1 merge790 (.A1(net518),
    .A2(net532),
    .A3(net652),
    .B1(net651),
    .X(net749));
 sky130_fd_sc_hd__a41o_1 merge791 (.A1(net242),
    .A2(net391),
    .A3(net388),
    .A4(net382),
    .B1(net961),
    .X(net750));
 sky130_fd_sc_hd__mux4_1 merge792 (.A0(net274),
    .A1(net968),
    .A2(net536),
    .A3(net539),
    .S0(net1064),
    .S1(net781),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 merge793 (.A0(net545),
    .A1(net1007),
    .A2(net1064),
    .A3(net398),
    .S0(net254),
    .S1(net1150),
    .X(net752));
 sky130_fd_sc_hd__mux4_1 merge794 (.A0(net382),
    .A1(net235),
    .A2(net1067),
    .A3(net258),
    .S0(net252),
    .S1(net1017),
    .X(net753));
 sky130_fd_sc_hd__a41o_1 merge795 (.A1(net643),
    .A2(net652),
    .A3(net642),
    .A4(net1121),
    .B1(net529),
    .X(net754));
 sky130_fd_sc_hd__mux4_1 merge796 (.A0(net249),
    .A1(net642),
    .A2(net522),
    .A3(net391),
    .S0(net549),
    .S1(net545),
    .X(net755));
 sky130_fd_sc_hd__a41o_1 merge797 (.A1(net513),
    .A2(net382),
    .A3(net107),
    .A4(net515),
    .B1(net391),
    .X(net756));
 sky130_fd_sc_hd__mux4_1 merge798 (.A0(net983),
    .A1(net380),
    .A2(net254),
    .A3(net543),
    .S0(net387),
    .S1(net547),
    .X(net757));
 sky130_fd_sc_hd__mux4_1 merge799 (.A0(net398),
    .A1(net396),
    .A2(net254),
    .A3(net518),
    .S0(net516),
    .S1(net519),
    .X(net758));
 sky130_fd_sc_hd__xnor2_1 merge800 (.A(net711),
    .B(net712),
    .Y(net759));
 sky130_fd_sc_hd__dfrbp_1 merge801 (.CLK(clknet_4_15_0_clk),
    .D(net678),
    .RESET_B(net661),
    .Q(net761),
    .Q_N(net760));
 sky130_fd_sc_hd__xnor2_1 merge802 (.A(net281),
    .B(net298),
    .Y(net762));
 sky130_fd_sc_hd__xnor2_1 merge803 (.A(net624),
    .B(net625),
    .Y(net763));
 sky130_fd_sc_hd__dfrbp_1 merge804 (.CLK(clknet_4_0_0_clk),
    .D(net215),
    .RESET_B(net216),
    .Q(net765),
    .Q_N(net764));
 sky130_fd_sc_hd__dfrtn_1 merge805 (.CLK_N(clknet_4_13_0_clk),
    .D(net753),
    .RESET_B(net392),
    .Q(net766));
 sky130_fd_sc_hd__xnor2_1 merge806 (.A(net602),
    .B(net606),
    .Y(net767));
 sky130_fd_sc_hd__dfrtp_2 merge807 (.CLK(clknet_4_15_0_clk),
    .D(net749),
    .RESET_B(net754),
    .Q(net768));
 sky130_fd_sc_hd__xnor2_1 merge808 (.A(net557),
    .B(net560),
    .Y(net769));
 sky130_fd_sc_hd__dfrtp_1 merge809 (.CLK(clknet_4_13_0_clk),
    .D(net751),
    .RESET_B(net752),
    .Q(net770));
 sky130_fd_sc_hd__xnor2_1 merge810 (.A(net347),
    .B(net353),
    .Y(net771));
 sky130_fd_sc_hd__xnor2_1 merge811 (.A(net578),
    .B(net582),
    .Y(net772));
 sky130_fd_sc_hd__xnor2_2 merge812 (.A(net493),
    .B(net497),
    .Y(net773));
 sky130_fd_sc_hd__xnor2_1 merge813 (.A(net684),
    .B(net686),
    .Y(net774));
 sky130_fd_sc_hd__dfrtp_2 merge814 (.CLK(clknet_4_13_0_clk),
    .D(net531),
    .RESET_B(net750),
    .Q(net775));
 sky130_fd_sc_hd__xnor2_1 merge815 (.A(net472),
    .B(net478),
    .Y(net776));
 sky130_fd_sc_hd__xnor2_1 merge816 (.A(net454),
    .B(net460),
    .Y(net777));
 sky130_fd_sc_hd__xnor2_1 merge817 (.A(net318),
    .B(net321),
    .Y(net778));
 sky130_fd_sc_hd__xnor2_1 merge818 (.A(net189),
    .B(net188),
    .Y(net779));
 sky130_fd_sc_hd__dfsbp_2 merge819 (.CLK(clknet_4_12_0_clk),
    .D(net423),
    .SET_B(net409),
    .Q(net781),
    .Q_N(net780));
 sky130_fd_sc_hd__dfsbp_2 merge820 (.CLK(clknet_4_5_0_clk),
    .SET_B(net251),
    .Q(net783),
    .Q_N(net253));
 sky130_fd_sc_hd__xnor2_1 merge821 (.A(net356),
    .B(net357),
    .Y(net784));
 sky130_fd_sc_hd__dfstp_2 merge822 (.CLK(clknet_4_4_0_clk),
    .D(net278),
    .SET_B(net264),
    .Q(net785));
 sky130_fd_sc_hd__dfstp_1 merge823 (.CLK(clknet_4_10_0_clk),
    .D(net732),
    .SET_B(net734),
    .Q(net786));
 sky130_fd_sc_hd__dfstp_1 merge824 (.CLK(clknet_4_1_0_clk),
    .D(net209),
    .SET_B(net204),
    .Q(net787));
 sky130_fd_sc_hd__xnor2_1 merge825 (.A(net431),
    .B(net425),
    .Y(net788));
 sky130_fd_sc_hd__xnor2_1 merge826 (.A(net746),
    .B(net610),
    .Y(net789));
 sky130_fd_sc_hd__xnor2_1 merge827 (.A(net367),
    .B(net322),
    .Y(net790));
 sky130_fd_sc_hd__xnor2_1 merge828 (.A(net566),
    .B(net599),
    .Y(net791));
 sky130_fd_sc_hd__dlrbn_1 merge829 (.D(net771),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net350),
    .Q_N(net792));
 sky130_fd_sc_hd__dlrbn_1 merge830 (.D(net218),
    .GATE_N(clknet_4_0_0_clk),
    .RESET_B(net219),
    .Q(net795),
    .Q_N(net794));
 sky130_fd_sc_hd__dlrbp_1 merge831 (.D(net755),
    .GATE(clknet_4_15_0_clk),
    .RESET_B(net681),
    .Q(net797),
    .Q_N(net796));
 sky130_fd_sc_hd__dlrbp_1 merge832 (.D(net439),
    .GATE(clknet_4_4_0_clk),
    .RESET_B(net305),
    .Q(net799),
    .Q_N(net798));
 sky130_fd_sc_hd__dlrtn_2 merge833 (.D(net757),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net677),
    .Q(net800));
 sky130_fd_sc_hd__dlrtn_1 merge834 (.D(net328),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net778),
    .Q(net801));
 sky130_fd_sc_hd__xnor2_4 merge835 (.A(net773),
    .B(net511),
    .Y(net802));
 sky130_fd_sc_hd__dlrtn_1 merge836 (.D(net464),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net467),
    .Q(net803));
 sky130_fd_sc_hd__xnor2_1 merge837 (.A(net687),
    .B(net705),
    .Y(net804));
 sky130_fd_sc_hd__xnor2_1 merge838 (.A(net698),
    .B(net577),
    .Y(net805));
 sky130_fd_sc_hd__xnor2_1 merge839 (.A(net592),
    .B(net727),
    .Y(net806));
 sky130_fd_sc_hd__dlrtp_1 merge840 (.D(net612),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net636),
    .Q(net1000));
 sky130_fd_sc_hd__xnor2_1 merge841 (.A(net735),
    .B(net634),
    .Y(net807));
 sky130_fd_sc_hd__dlrtp_1 merge842 (.D(net360),
    .GATE(clknet_4_0_0_clk),
    .RESET_B(net364),
    .Q(net808));
 sky130_fd_sc_hd__xnor2_1 merge843 (.A(net485),
    .B(net483),
    .Y(net809));
 sky130_fd_sc_hd__xnor2_1 merge844 (.A(net571),
    .B(net621),
    .Y(net810));
 sky130_fd_sc_hd__xnor2_1 merge845 (.A(net572),
    .B(net725),
    .Y(net811));
 sky130_fd_sc_hd__dlrtp_2 merge846 (.D(net421),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net424),
    .Q(net812));
 sky130_fd_sc_hd__xnor2_1 merge847 (.A(net716),
    .B(net631),
    .Y(net813));
 sky130_fd_sc_hd__xnor2_1 merge848 (.A(net482),
    .B(net507),
    .Y(net814));
 sky130_fd_sc_hd__edfxbp_1 merge849 (.CLK(clknet_4_13_0_clk),
    .D(net756),
    .DE(net758),
    .Q(net816),
    .Q_N(net815));
 sky130_fd_sc_hd__edfxtp_1 merge850 (.CLK(clknet_4_11_0_clk),
    .D(net576),
    .DE(net810),
    .Q(net817));
 sky130_fd_sc_hd__xnor2_1 merge851 (.A(net737),
    .B(net722),
    .Y(net818));
 sky130_fd_sc_hd__sdlclkp_1 merge852 (.CLK(clknet_4_4_0_clk),
    .GATE(net146),
    .SCE(net180),
    .GCLK(net819));
 sky130_fd_sc_hd__xnor2_1 merge853 (.A(net584),
    .B(net614),
    .Y(net820));
 sky130_fd_sc_hd__xnor2_1 merge854 (.A(net300),
    .B(net304),
    .Y(net821));
 sky130_fd_sc_hd__sdlclkp_2 merge855 (.CLK(clknet_4_8_0_clk),
    .GATE(net616),
    .SCE(net627),
    .GCLK(net822));
 sky130_fd_sc_hd__sdlclkp_4 merge856 (.CLK(clknet_4_0_0_clk),
    .GATE(net220),
    .SCE(net227),
    .GCLK(net823));
 sky130_fd_sc_hd__xnor2_1 merge857 (.A(net745),
    .B(net589),
    .Y(net824));
 sky130_fd_sc_hd__dfrbp_2 merge858 (.CLK(clknet_4_1_0_clk),
    .D(net187),
    .RESET_B(net779),
    .Q(net826),
    .Q_N(net825));
 sky130_fd_sc_hd__dfrbp_2 merge859 (.CLK(clknet_4_4_0_clk),
    .D(net271),
    .RESET_B(net276),
    .Q(net828),
    .Q_N(net827));
 sky130_fd_sc_hd__dfrtn_1 merge860 (.CLK_N(clknet_4_0_0_clk),
    .D(net332),
    .RESET_B(net790),
    .Q(net829));
 sky130_fd_sc_hd__xnor2_1 merge861 (.A(net618),
    .B(net506),
    .Y(net830));
 sky130_fd_sc_hd__dfrtp_4 merge862 (.CLK(clknet_4_15_0_clk),
    .D(net813),
    .RESET_B(net664),
    .Q(net831));
 sky130_fd_sc_hd__dfrtp_4 merge863 (.CLK(clknet_4_11_0_clk),
    .D(net811),
    .RESET_B(net791),
    .Q(net832));
 sky130_fd_sc_hd__xnor2_1 merge864 (.A(net736),
    .B(net505),
    .Y(net833));
 sky130_fd_sc_hd__dfrtp_1 merge865 (.CLK(clknet_4_2_0_clk),
    .D(net503),
    .RESET_B(net337),
    .Q(net834));
 sky130_fd_sc_hd__dfsbp_1 merge866 (.CLK(clknet_4_6_0_clk),
    .D(net457),
    .SET_B(net777),
    .Q(net836),
    .Q_N(net835));
 sky130_fd_sc_hd__dfsbp_1 merge867 (.CLK(clknet_4_14_0_clk),
    .D(net672),
    .SET_B(net804),
    .Q(net838),
    .Q_N(net837));
 sky130_fd_sc_hd__xnor2_1 merge868 (.A(net747),
    .B(net740),
    .Y(net839));
 sky130_fd_sc_hd__dfstp_1 merge869 (.CLK(clknet_4_15_0_clk),
    .D(net697),
    .SET_B(net774),
    .Q(net840));
 sky130_fd_sc_hd__dfstp_1 merge870 (.CLK(clknet_4_8_0_clk),
    .D(net579),
    .SET_B(net632),
    .Q(net841));
 sky130_fd_sc_hd__dfstp_2 merge871 (.CLK(clknet_4_7_0_clk),
    .D(net330),
    .SET_B(net290),
    .Q(net842));
 sky130_fd_sc_hd__dlrbn_1 merge872 (.D(net805),
    .GATE_N(clknet_4_11_0_clk),
    .RESET_B(net759),
    .Q(net843),
    .Q_N(net986));
 sky130_fd_sc_hd__dlrbn_1 merge873 (.D(net488),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net630),
    .Q(net845),
    .Q_N(net844));
 sky130_fd_sc_hd__dlrbp_1 merge874 (.D(net689),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net802),
    .Q(net846),
    .Q_N(net1006));
 sky130_fd_sc_hd__dlrbp_1 merge875 (.D(net809),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net502),
    .Q(net848),
    .Q_N(net847));
 sky130_fd_sc_hd__dlrtn_2 merge876 (.D(net690),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net833),
    .Q(net849));
 sky130_fd_sc_hd__dlrtn_1 merge877 (.D(net615),
    .GATE_N(clknet_4_8_0_clk),
    .RESET_B(net480),
    .Q(net850));
 sky130_fd_sc_hd__dlrtn_1 merge878 (.D(net348),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net494),
    .Q(net851));
 sky130_fd_sc_hd__dlrtp_2 merge879 (.D(net704),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net688),
    .Q(net852));
 sky130_fd_sc_hd__dlrtp_1 merge880 (.D(net474),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net824),
    .Q(net853));
 sky130_fd_sc_hd__dlrtp_1 merge881 (.D(net788),
    .GATE(clknet_4_7_0_clk),
    .RESET_B(net435),
    .Q(net854));
 sky130_fd_sc_hd__edfxbp_1 merge882 (.CLK(clknet_4_8_0_clk),
    .D(net763),
    .DE(net767),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__edfxtp_1 merge883 (.CLK(clknet_4_0_0_clk),
    .D(net228),
    .DE(net784),
    .Q(net857));
 sky130_fd_sc_hd__sdlclkp_1 merge884 (.CLK(clknet_4_11_0_clk),
    .GATE(net593),
    .SCE(net806),
    .GCLK(net858));
 sky130_fd_sc_hd__sdlclkp_2 merge885 (.CLK(clknet_4_7_0_clk),
    .GATE(net762),
    .SCE(net821),
    .GCLK(net859));
 sky130_fd_sc_hd__sdlclkp_4 merge886 (.CLK(clknet_4_10_0_clk),
    .GATE(net830),
    .SCE(net818),
    .GCLK(net994));
 sky130_fd_sc_hd__dfrbp_1 merge887 (.CLK(clknet_4_11_0_clk),
    .D(net691),
    .RESET_B(net820),
    .Q(net861),
    .Q_N(net860));
 sky130_fd_sc_hd__dfrbp_1 merge888 (.CLK(clknet_4_9_0_clk),
    .D(net772),
    .RESET_B(net769),
    .Q(net863),
    .Q_N(net862));
 sky130_fd_sc_hd__dfrtn_1 merge889 (.CLK_N(clknet_4_3_0_clk),
    .D(net776),
    .RESET_B(net491),
    .Q(net864));
 sky130_fd_sc_hd__dfrtp_4 merge890 (.CLK(clknet_4_10_0_clk),
    .D(net789),
    .RESET_B(net674),
    .Q(net865));
 sky130_fd_sc_hd__dfrtp_4 merge891 (.CLK(clknet_4_3_0_clk),
    .D(net814),
    .RESET_B(net449),
    .Q(net866));
 sky130_fd_sc_hd__dfrtp_1 merge892 (.CLK(clknet_4_2_0_clk),
    .RESET_B(net373),
    .Q(net375));
 sky130_fd_sc_hd__dfsbp_1 merge893 (.CLK(clknet_4_8_0_clk),
    .D(net613),
    .SET_B(net601),
    .Q(net869),
    .Q_N(net868));
 sky130_fd_sc_hd__dfsbp_1 merge894 (.CLK(clknet_4_10_0_clk),
    .D(net839),
    .SET_B(net807),
    .Q(net871),
    .Q_N(net870));
 sky130_fd_sc_hd__dfstp_2 merge895 (.CLK(clknet_4_3_0_clk),
    .D(net349),
    .SET_B(net343),
    .Q(net872));
 sky130_fd_sc_hd__dfxbp_1 s896 (.CLK(clknet_4_0_0_clk),
    .D(net101),
    .Q(net874),
    .Q_N(net873));
 sky130_fd_sc_hd__dfxbp_1 s897 (.CLK(clknet_4_0_0_clk),
    .D(net211),
    .Q(net876),
    .Q_N(net875));
 sky130_fd_sc_hd__dfxtp_1 s898 (.CLK(clknet_4_0_0_clk),
    .D(net223),
    .Q(net877));
 sky130_fd_sc_hd__dfxtp_2 s899 (.CLK(clknet_4_5_0_clk),
    .D(net277),
    .Q(net878));
 sky130_fd_sc_hd__dfxtp_1 s900 (.CLK(clknet_4_5_0_clk),
    .D(net279),
    .Q(net879));
 sky130_fd_sc_hd__dlclkp_1 s901 (.CLK(clknet_4_5_0_clk),
    .GATE(net282),
    .GCLK(net880));
 sky130_fd_sc_hd__dlclkp_2 s902 (.CLK(clknet_4_4_0_clk),
    .GATE(net299),
    .GCLK(net881));
 sky130_fd_sc_hd__dlclkp_4 s903 (.CLK(clknet_4_7_0_clk),
    .GATE(net303),
    .GCLK(net882));
 sky130_fd_sc_hd__dlxbn_1 s904 (.D(net314),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net884),
    .Q_N(net883));
 sky130_fd_sc_hd__dlxbn_2 s905 (.D(net319),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net886),
    .Q_N(net885));
 sky130_fd_sc_hd__dlxbp_1 s906 (.D(net325),
    .GATE(clknet_4_9_0_clk),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__dlxtn_1 s907 (.D(net326),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net889));
 sky130_fd_sc_hd__dlxtn_1 s908 (.D(net329),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net890));
 sky130_fd_sc_hd__dlxtn_1 s909 (.D(net340),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net891));
 sky130_fd_sc_hd__dlxtp_1 s910 (.D(net342),
    .GATE(clknet_4_3_0_clk),
    .Q(net892));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s911 (.D(net368),
    .SLEEP_B(clknet_4_2_0_clk),
    .Q(net893));
 sky130_fd_sc_hd__dfxbp_1 s912 (.CLK(clknet_4_2_0_clk),
    .D(net369),
    .Q(net895),
    .Q_N(net894));
 sky130_fd_sc_hd__dfxbp_1 s913 (.CLK(clknet_4_2_0_clk),
    .D(net370),
    .Q(net897),
    .Q_N(net896));
 sky130_fd_sc_hd__dfxtp_1 s914 (.CLK(clknet_4_2_0_clk),
    .D(net372),
    .Q(net898));
 sky130_fd_sc_hd__dfxtp_2 s915 (.CLK(clknet_4_12_0_clk),
    .D(net428),
    .Q(net899));
 sky130_fd_sc_hd__dfxtp_1 s916 (.CLK(clknet_4_12_0_clk),
    .D(net444),
    .Q(net900));
 sky130_fd_sc_hd__dlclkp_1 s917 (.CLK(clknet_4_12_0_clk),
    .GATE(net445),
    .GCLK(net901));
 sky130_fd_sc_hd__dlclkp_2 s918 (.CLK(clknet_4_6_0_clk),
    .GATE(net450),
    .GCLK(net902));
 sky130_fd_sc_hd__dlclkp_4 s919 (.CLK(clknet_4_9_0_clk),
    .GATE(net451),
    .GCLK(net903));
 sky130_fd_sc_hd__dlxbn_2 s920 (.D(net459),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net905),
    .Q_N(net904));
 sky130_fd_sc_hd__dlxbn_2 s921 (.D(net461),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net907),
    .Q_N(net906));
 sky130_fd_sc_hd__dlxbp_1 s922 (.D(net462),
    .GATE(clknet_4_9_0_clk),
    .Q(net909),
    .Q_N(net908));
 sky130_fd_sc_hd__dlxtn_1 s923 (.D(net471),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net910));
 sky130_fd_sc_hd__dlxtn_1 s924 (.D(net479),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net911));
 sky130_fd_sc_hd__dlxtn_1 s925 (.D(net484),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net912));
 sky130_fd_sc_hd__dlxtp_1 s926 (.D(net486),
    .GATE(clknet_4_3_0_clk),
    .Q(net913));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s927 (.D(net490),
    .SLEEP_B(clknet_4_3_0_clk),
    .Q(net914));
 sky130_fd_sc_hd__dfxbp_1 s928 (.CLK(clknet_4_2_0_clk),
    .D(net498),
    .Q(net916),
    .Q_N(net915));
 sky130_fd_sc_hd__dfxbp_1 s929 (.CLK(clknet_4_2_0_clk),
    .D(net501),
    .Q(net918),
    .Q_N(net917));
 sky130_fd_sc_hd__dfxtp_1 s930 (.CLK(clknet_4_13_0_clk),
    .D(net512),
    .Q(net919));
 sky130_fd_sc_hd__dfxtp_1 s931 (.CLK(clknet_4_13_0_clk),
    .D(net548),
    .Q(net920));
 sky130_fd_sc_hd__dfxtp_1 s932 (.CLK(clknet_4_13_0_clk),
    .D(net550),
    .Q(net921));
 sky130_fd_sc_hd__dlclkp_1 s933 (.CLK(clknet_4_12_0_clk),
    .GATE(net564),
    .GCLK(net922));
 sky130_fd_sc_hd__dlclkp_2 s934 (.CLK(clknet_4_14_0_clk),
    .GATE(net565),
    .GCLK(net923));
 sky130_fd_sc_hd__dlclkp_4 s935 (.CLK(clknet_4_14_0_clk),
    .GATE(net569),
    .GCLK(net924));
 sky130_fd_sc_hd__dlxbn_1 s936 (.D(net573),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net926),
    .Q_N(net925));
 sky130_fd_sc_hd__dlxbn_1 s937 (.D(net575),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net991),
    .Q_N(net927));
 sky130_fd_sc_hd__dlxbp_1 s938 (.D(net580),
    .GATE(clknet_4_9_0_clk),
    .Q(net929),
    .Q_N(net928));
 sky130_fd_sc_hd__dlxtn_4 s939 (.D(net581),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net930));
 sky130_fd_sc_hd__dlxtn_1 s940 (.D(net585),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net931));
 sky130_fd_sc_hd__dlxtn_1 s941 (.D(net586),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net932));
 sky130_fd_sc_hd__dlxtp_1 s942 (.D(net587),
    .GATE(clknet_4_11_0_clk),
    .Q(net933));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s943 (.D(net590),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net934));
 sky130_fd_sc_hd__dfxbp_1 s944 (.CLK(clknet_4_10_0_clk),
    .D(net591),
    .Q(net936),
    .Q_N(net935));
 sky130_fd_sc_hd__dfxbp_1 s945 (.CLK(clknet_4_8_0_clk),
    .D(net598),
    .Q(net938),
    .Q_N(net937));
 sky130_fd_sc_hd__dfxtp_1 s946 (.CLK(clknet_4_8_0_clk),
    .D(net626),
    .Q(net939));
 sky130_fd_sc_hd__dfxtp_1 s947 (.CLK(clknet_4_15_0_clk),
    .D(net658),
    .Q(net940));
 sky130_fd_sc_hd__dfxtp_1 s948 (.CLK(clknet_4_15_0_clk),
    .D(net669),
    .Q(net941));
 sky130_fd_sc_hd__dlclkp_1 s949 (.CLK(clknet_4_14_0_clk),
    .GATE(net685),
    .GCLK(net942));
 sky130_fd_sc_hd__dlclkp_2 s950 (.CLK(clknet_4_14_0_clk),
    .GATE(net692),
    .GCLK(net943));
 sky130_fd_sc_hd__dlclkp_4 s951 (.CLK(clknet_4_14_0_clk),
    .GATE(net695),
    .GCLK(net944));
 sky130_fd_sc_hd__dlxbn_1 s952 (.D(net699),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net946),
    .Q_N(net945));
 sky130_fd_sc_hd__dlxbn_1 s953 (.D(net701),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net948),
    .Q_N(net947));
 sky130_fd_sc_hd__dlxbp_1 s954 (.D(net702),
    .GATE(clknet_4_14_0_clk),
    .Q(net950),
    .Q_N(net949));
 sky130_fd_sc_hd__dlxtn_1 s955 (.D(net707),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net951));
 sky130_fd_sc_hd__dlxtn_2 s956 (.D(net714),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net952));
 sky130_fd_sc_hd__dlxtn_1 s957 (.D(net717),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net953));
 sky130_fd_sc_hd__dlxtp_1 s958 (.D(net720),
    .GATE(clknet_4_11_0_clk),
    .Q(net954));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s959 (.D(net724),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net955));
 sky130_fd_sc_hd__dfxbp_1 s960 (.CLK(clknet_4_10_0_clk),
    .D(net729),
    .Q(net957),
    .Q_N(net956));
 sky130_fd_sc_hd__dfxbp_1 s961 (.CLK(clknet_4_10_0_clk),
    .D(net741),
    .Q(net959),
    .Q_N(net958));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(in0),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1),
    .X(net961));
 sky130_fd_sc_hd__buf_1 input3 (.A(in10),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in11),
    .X(net963));
 sky130_fd_sc_hd__buf_8 input5 (.A(in12),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(in13),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in15),
    .X(net967));
 sky130_fd_sc_hd__buf_8 input9 (.A(in16),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(in17),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in18),
    .X(net970));
 sky130_fd_sc_hd__buf_2 input12 (.A(in19),
    .X(net971));
 sky130_fd_sc_hd__buf_12 input13 (.A(in2),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in20),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in21),
    .X(net974));
 sky130_fd_sc_hd__buf_6 input16 (.A(in22),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_8 input17 (.A(in23),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_8 input18 (.A(in24),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(in3),
    .X(net978));
 sky130_fd_sc_hd__buf_8 input20 (.A(in4),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in5),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in6),
    .X(net981));
 sky130_fd_sc_hd__buf_6 input23 (.A(in7),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in8),
    .X(net983));
 sky130_fd_sc_hd__buf_4 input25 (.A(in9),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(clknet_1_0__leaf_net985),
    .X(out0));
 sky130_fd_sc_hd__buf_2 output27 (.A(net986),
    .X(out1));
 sky130_fd_sc_hd__buf_2 output28 (.A(net987),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output29 (.A(net988),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output30 (.A(net1066),
    .X(out13));
 sky130_fd_sc_hd__buf_2 output31 (.A(net1052),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output32 (.A(net991),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output33 (.A(net992),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output34 (.A(net993),
    .X(out18));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(clknet_1_0__leaf_net994),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output36 (.A(net995),
    .X(out2));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(clknet_1_0__leaf_net996),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net997),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output39 (.A(net998),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output40 (.A(net999),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output41 (.A(net1000),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output42 (.A(net1001),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output43 (.A(net1002),
    .X(out5));
 sky130_fd_sc_hd__buf_2 output44 (.A(net1065),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output45 (.A(net1004),
    .X(out7));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net1005),
    .X(out8));
 sky130_fd_sc_hd__buf_2 output47 (.A(net1006),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net520),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout49 (.A(net422),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net395),
    .X(net1009));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net270),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net270),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout53 (.A(net246),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net556),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net283),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 max_cap56 (.A(net245),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 max_cap57 (.A(net379),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net1019),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net261),
    .X(net1019));
 sky130_fd_sc_hd__buf_8 fanout61 (.A(net123),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 max_cap62 (.A(net84),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 max_cap63 (.A(net242),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net169),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net160),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net160),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net1116),
    .X(net1026));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net119),
    .X(net1027));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net119),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(net81),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net55),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_8 fanout73 (.A(net238),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 max_cap74 (.A(net131),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net66),
    .X(net1034));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(net34),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 max_cap77 (.A(net988),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net33),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(net33),
    .X(net1038));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(net116),
    .X(net1039));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net116),
    .X(net1040));
 sky130_fd_sc_hd__buf_6 fanout82 (.A(net50),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_8 fanout83 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(net115),
    .X(net1043));
 sky130_fd_sc_hd__buf_12 fanout85 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net112),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 max_cap87 (.A(net40),
    .X(net1046));
 sky130_fd_sc_hd__buf_6 fanout88 (.A(net24),
    .X(net1047));
 sky130_fd_sc_hd__buf_4 max_cap89 (.A(net993),
    .X(net1048));
 sky130_fd_sc_hd__buf_4 max_cap90 (.A(net21),
    .X(net1049));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(net153),
    .X(net1050));
 sky130_fd_sc_hd__buf_4 max_cap92 (.A(net39),
    .X(net1051));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(net990),
    .X(net1053));
 sky130_fd_sc_hd__buf_12 fanout95 (.A(net109),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 wire96 (.A(net19),
    .X(net1055));
 sky130_fd_sc_hd__buf_4 max_cap97 (.A(net14),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net147),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 max_cap99 (.A(net22),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net385),
    .X(net1059));
 sky130_fd_sc_hd__buf_4 max_cap101 (.A(net7),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 wire102 (.A(net3),
    .X(net1061));
 sky130_fd_sc_hd__buf_4 max_cap103 (.A(net2),
    .X(net1062));
 sky130_fd_sc_hd__buf_8 max_cap104 (.A(net107),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__buf_4 fanout106 (.A(net1003),
    .X(net1065));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net989),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net1070),
    .X(net1067));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net1070),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net381),
    .X(net1070));
 sky130_fd_sc_hd__buf_4 max_cap112 (.A(net12),
    .X(net1071));
 sky130_fd_sc_hd__buf_4 max_cap113 (.A(net10),
    .X(net1072));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net6),
    .X(net1073));
 sky130_fd_sc_hd__buf_4 max_cap115 (.A(net236),
    .X(net1074));
 sky130_fd_sc_hd__buf_12 max_cap116 (.A(net104),
    .X(net1075));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net879),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net879),
    .X(net1077));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net878),
    .X(net1078));
 sky130_fd_sc_hd__buf_4 max_cap120 (.A(net766),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net408),
    .X(net1080));
 sky130_fd_sc_hd__buf_4 max_cap122 (.A(net8),
    .X(net1081));
 sky130_fd_sc_hd__buf_4 max_cap123 (.A(net1083),
    .X(net1082));
 sky130_fd_sc_hd__buf_4 max_cap124 (.A(net5),
    .X(net1083));
 sky130_fd_sc_hd__buf_4 max_cap125 (.A(net4),
    .X(net1084));
 sky130_fd_sc_hd__buf_4 max_cap126 (.A(net0),
    .X(net1085));
 sky130_fd_sc_hd__buf_4 max_cap127 (.A(net105),
    .X(net1086));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net102),
    .X(net1087));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(net967),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net966),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(net963),
    .X(net1091));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net1093),
    .X(net1092));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net962),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_8 fanout135 (.A(net984),
    .X(net1094));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(net983),
    .X(net1095));
 sky130_fd_sc_hd__buf_12 fanout137 (.A(net982),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net981),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_8 fanout139 (.A(net980),
    .X(net1098));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(net961),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_8 fanout141 (.A(net978),
    .X(net1100));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net974),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net974),
    .X(net1102));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net973),
    .X(net1103));
 sky130_fd_sc_hd__buf_12 fanout145 (.A(net972),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(net971),
    .X(net1105));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net970),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(net960),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net944 (.A(net944),
    .X(clknet_0_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_0__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_1__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net696 (.A(net696),
    .X(clknet_0_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_0__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net696 (.A(clknet_0_net696),
    .X(clknet_1_1__leaf_net696));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net709 (.A(net709),
    .X(clknet_0_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_0__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net709 (.A(clknet_0_net709),
    .X(clknet_1_1__leaf_net709));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net858 (.A(net858),
    .X(clknet_0_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_0__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net858 (.A(clknet_0_net858),
    .X(clknet_1_1__leaf_net858));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net597 (.A(net597),
    .X(clknet_0_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_0__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net597 (.A(clknet_0_net597),
    .X(clknet_1_1__leaf_net597));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net611 (.A(net611),
    .X(clknet_0_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_0__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net611 (.A(clknet_0_net611),
    .X(clknet_1_1__leaf_net611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net822 (.A(net822),
    .X(clknet_0_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_0__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net822 (.A(clknet_0_net822),
    .X(clknet_1_1__leaf_net822));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net994 (.A(net994),
    .X(clknet_0_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_0__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net994 (.A(clknet_0_net994),
    .X(clknet_1_1__leaf_net994));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net595 (.A(net595),
    .X(clknet_0_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_0__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net595 (.A(clknet_0_net595),
    .X(clknet_1_1__leaf_net595));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net607 (.A(net607),
    .X(clknet_0_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net607 (.A(clknet_0_net607),
    .X(clknet_1_0__leaf_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net607 (.A(clknet_0_net607),
    .X(clknet_1_1__leaf_net607));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net943 (.A(net943),
    .X(clknet_0_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net943 (.A(clknet_0_net943),
    .X(clknet_1_0__leaf_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net943 (.A(clknet_0_net943),
    .X(clknet_1_1__leaf_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net703 (.A(net703),
    .X(clknet_0_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_0__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net703 (.A(clknet_0_net703),
    .X(clknet_1_1__leaf_net703));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net942 (.A(net942),
    .X(clknet_0_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_0__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_1__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net570 (.A(net570),
    .X(clknet_0_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_0__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net570 (.A(clknet_0_net570),
    .X(clknet_1_1__leaf_net570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net923 (.A(net923),
    .X(clknet_0_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net903 (.A(net903),
    .X(clknet_0_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net903 (.A(clknet_0_net903),
    .X(clknet_1_0__leaf_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net903 (.A(clknet_0_net903),
    .X(clknet_1_1__leaf_net903));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net902 (.A(net902),
    .X(clknet_0_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_0__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net902 (.A(clknet_0_net902),
    .X(clknet_1_1__leaf_net902));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net596 (.A(net596),
    .X(clknet_0_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_0__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net596 (.A(clknet_0_net596),
    .X(clknet_1_1__leaf_net596));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net706 (.A(net706),
    .X(clknet_0_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_0__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net706 (.A(clknet_0_net706),
    .X(clknet_1_1__leaf_net706));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net562 (.A(net562),
    .X(clknet_0_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_0__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net562 (.A(clknet_0_net562),
    .X(clknet_1_1__leaf_net562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net567 (.A(net567),
    .X(clknet_0_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_0__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net567 (.A(clknet_0_net567),
    .X(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net693 (.A(net693),
    .X(clknet_0_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_0__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net693 (.A(clknet_0_net693),
    .X(clknet_1_1__leaf_net693));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net561 (.A(net561),
    .X(clknet_0_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_0__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net561 (.A(clknet_0_net561),
    .X(clknet_1_1__leaf_net561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net882 (.A(net882),
    .X(clknet_0_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net882 (.A(clknet_0_net882),
    .X(clknet_1_1__leaf_net882));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net700 (.A(net700),
    .X(clknet_0_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_0__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net700 (.A(clknet_0_net700),
    .X(clknet_1_1__leaf_net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net859 (.A(net859),
    .X(clknet_0_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_0__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net859 (.A(clknet_0_net859),
    .X(clknet_1_1__leaf_net859));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net436 (.A(net436),
    .X(clknet_0_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_0__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net436 (.A(clknet_0_net436),
    .X(clknet_1_1__leaf_net436));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net327 (.A(net327),
    .X(clknet_0_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_0__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net327 (.A(clknet_0_net327),
    .X(clknet_1_1__leaf_net327));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net313 (.A(net313),
    .X(clknet_0_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_0__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net313 (.A(clknet_0_net313),
    .X(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net297 (.A(net297),
    .X(clknet_0_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_0__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net297 (.A(clknet_0_net297),
    .X(clknet_1_1__leaf_net297));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net881 (.A(net881),
    .X(clknet_0_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net881 (.A(clknet_0_net881),
    .X(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net881 (.A(clknet_0_net881),
    .X(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net455 (.A(net455),
    .X(clknet_0_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_0__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net455 (.A(clknet_0_net455),
    .X(clknet_1_1__leaf_net455));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net985 (.A(net985),
    .X(clknet_0_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_0__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net985 (.A(clknet_0_net985),
    .X(clknet_1_1__leaf_net985));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net286 (.A(net286),
    .X(clknet_0_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_0__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net286 (.A(clknet_0_net286),
    .X(clknet_1_1__leaf_net286));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net880 (.A(net880),
    .X(clknet_0_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_0__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net880 (.A(clknet_0_net880),
    .X(clknet_1_1__leaf_net880));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net339 (.A(net339),
    .X(clknet_0_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_0__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net339 (.A(clknet_0_net339),
    .X(clknet_1_1__leaf_net339));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net296 (.A(net296),
    .X(clknet_0_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_0__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net296 (.A(clknet_0_net296),
    .X(clknet_1_1__leaf_net296));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net823 (.A(net823),
    .X(clknet_0_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_0__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net823 (.A(clknet_0_net823),
    .X(clknet_1_1__leaf_net823));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net234 (.A(net234),
    .X(clknet_0_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_0__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net234 (.A(clknet_0_net234),
    .X(clknet_1_1__leaf_net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net225 (.A(net225),
    .X(clknet_0_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_0__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net225 (.A(clknet_0_net225),
    .X(clknet_1_1__leaf_net225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net222 (.A(net222),
    .X(clknet_0_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_0__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net222 (.A(clknet_0_net222),
    .X(clknet_1_1__leaf_net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net499 (.A(net499),
    .X(clknet_0_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_0__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net499 (.A(clknet_0_net499),
    .X(clknet_1_1__leaf_net499));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net231 (.A(net231),
    .X(clknet_0_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_0__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net231 (.A(clknet_0_net231),
    .X(clknet_1_1__leaf_net231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net226 (.A(net226),
    .X(clknet_0_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_0__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net226 (.A(clknet_0_net226),
    .X(clknet_1_1__leaf_net226));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net233 (.A(net233),
    .X(clknet_0_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_0__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net233 (.A(clknet_0_net233),
    .X(clknet_1_1__leaf_net233));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net819 (.A(net819),
    .X(clknet_0_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_0__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_1__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net331 (.A(net331),
    .X(clknet_0_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_0__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net331 (.A(clknet_0_net331),
    .X(clknet_1_1__leaf_net331));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net635 (.A(net635),
    .X(clknet_0_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_0__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net635 (.A(clknet_0_net635),
    .X(clknet_1_1__leaf_net635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net996 (.A(net996),
    .X(clknet_0_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net996 (.A(clknet_0_net996),
    .X(clknet_1_0__leaf_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net996 (.A(clknet_0_net996),
    .X(clknet_1_1__leaf_net996));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net352 (.A(net352),
    .X(clknet_0_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_0__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net352 (.A(clknet_0_net352),
    .X(clknet_1_1__leaf_net352));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net496 (.A(net496),
    .X(clknet_0_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_0__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net496 (.A(clknet_0_net496),
    .X(clknet_1_1__leaf_net496));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net309 (.A(net309),
    .X(clknet_0_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_0__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net309 (.A(clknet_0_net309),
    .X(clknet_1_1__leaf_net309));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net289 (.A(net289),
    .X(clknet_0_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_0__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net289 (.A(clknet_0_net289),
    .X(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net489 (.A(net489),
    .X(clknet_0_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_0__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net489 (.A(clknet_0_net489),
    .X(clknet_1_1__leaf_net489));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net609 (.A(net609),
    .X(clknet_0_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_0__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net609 (.A(clknet_0_net609),
    .X(clknet_1_1__leaf_net609));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net605 (.A(net605),
    .X(clknet_0_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_0__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net605 (.A(clknet_0_net605),
    .X(clknet_1_1__leaf_net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net604 (.A(net604),
    .X(clknet_0_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_0__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net604 (.A(clknet_0_net604),
    .X(clknet_1_1__leaf_net604));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net470 (.A(net470),
    .X(clknet_0_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net470 (.A(net1145),
    .X(clknet_1_0__leaf_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net470 (.A(clknet_0_net470),
    .X(clknet_1_1__leaf_net470));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net500 (.A(net500),
    .X(clknet_0_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_0__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net500 (.A(clknet_0_net500),
    .X(clknet_1_1__leaf_net500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net504 (.A(net504),
    .X(clknet_0_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_0__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net504 (.A(clknet_0_net504),
    .X(clknet_1_1__leaf_net504));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net469 (.A(net469),
    .X(clknet_0_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_0__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net469 (.A(clknet_0_net469),
    .X(clknet_1_1__leaf_net469));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net442 (.A(net442),
    .X(clknet_0_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_0__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net442 (.A(clknet_0_net442),
    .X(clknet_1_1__leaf_net442));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net447 (.A(net447),
    .X(clknet_0_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_0__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net447 (.A(clknet_0_net447),
    .X(clknet_1_1__leaf_net447));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net163 (.A(net163),
    .X(clknet_0_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_0__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net163 (.A(clknet_0_net163),
    .X(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net317 (.A(net317),
    .X(clknet_0_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_0__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net317 (.A(clknet_0_net317),
    .X(clknet_1_1__leaf_net317));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net315 (.A(net315),
    .X(clknet_0_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_0__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net315 (.A(clknet_0_net315),
    .X(clknet_1_1__leaf_net315));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net221 (.A(net221),
    .X(clknet_0_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_0__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net221 (.A(clknet_0_net221),
    .X(clknet_1_1__leaf_net221));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net192 (.A(net192),
    .X(clknet_0_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_0__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net192 (.A(clknet_0_net192),
    .X(clknet_1_1__leaf_net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net174 (.A(net174),
    .X(clknet_0_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net174 (.A(clknet_0_net174),
    .X(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net456 (.A(net456),
    .X(clknet_0_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_0__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net456 (.A(clknet_0_net456),
    .X(clknet_1_1__leaf_net456));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net320 (.A(net320),
    .X(clknet_0_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_0__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net320 (.A(clknet_0_net320),
    .X(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net186 (.A(net186),
    .X(clknet_0_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_0__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net186 (.A(clknet_0_net186),
    .X(clknet_1_1__leaf_net186));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net185 (.A(net185),
    .X(clknet_0_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_0__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net185 (.A(clknet_0_net185),
    .X(clknet_1_1__leaf_net185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net181 (.A(net181),
    .X(clknet_0_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_0__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net181 (.A(clknet_0_net181),
    .X(clknet_1_1__leaf_net181));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net175 (.A(net175),
    .X(clknet_0_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_0__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net175 (.A(clknet_0_net175),
    .X(clknet_1_1__leaf_net175));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net152 (.A(net152),
    .X(clknet_0_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_0__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net152 (.A(clknet_0_net152),
    .X(clknet_1_1__leaf_net152));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net167 (.A(net167),
    .X(clknet_0_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_0__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net167 (.A(clknet_0_net167),
    .X(clknet_1_1__leaf_net167));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net177 (.A(net177),
    .X(clknet_0_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net177 (.A(clknet_0_net177),
    .X(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net600 (.A(net600),
    .X(clknet_0_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_0__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net600 (.A(clknet_0_net600),
    .X(clknet_1_1__leaf_net600));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net351 (.A(net351),
    .X(clknet_0_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_0__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net351 (.A(clknet_0_net351),
    .X(clknet_1_1__leaf_net351));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net182 (.A(net182),
    .X(clknet_0_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_0__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net182 (.A(clknet_0_net182),
    .X(clknet_1_1__leaf_net182));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net179 (.A(net179),
    .X(clknet_0_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_0__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net179 (.A(clknet_0_net179),
    .X(clknet_1_1__leaf_net179));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net165 (.A(net165),
    .X(clknet_0_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net165 (.A(clknet_0_net165),
    .X(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net191 (.A(net191),
    .X(clknet_0_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_0__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net191 (.A(clknet_0_net191),
    .X(clknet_1_1__leaf_net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net203 (.A(net203),
    .X(clknet_0_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net203 (.A(clknet_0_net203),
    .X(clknet_1_1__leaf_net203));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net161 (.A(net161),
    .X(clknet_0_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net161 (.A(clknet_0_net161),
    .X(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net437 (.A(net437),
    .X(clknet_0_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_0__leaf_net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net437 (.A(clknet_0_net437),
    .X(clknet_1_1__leaf_net437));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net121),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net1108),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net1108),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net1179),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net1111),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net1112),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net123),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1114),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net119),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1182),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net1182),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net104),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1119),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1119),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net1130),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net108),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net108),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net122),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net1125),
    .X(net1126));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer20 (.A(net1185),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net1127),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net1128),
    .X(net1129));
 sky130_fd_sc_hd__a21bo_1 clone23 (.A1(net1144),
    .A2(net1096),
    .B1_N(net1165),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net111),
    .X(net1131));
 sky130_fd_sc_hd__buf_12 rebuffer25 (.A(net1143),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net113),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net1133),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net1134),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net1135),
    .X(net1136));
 sky130_fd_sc_hd__clkbuf_1 clone30 (.A(net119),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_1 clone31 (.A(net109),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_4 clone32 (.A(net982),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(net1020),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net1140),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net117),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(net1142),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_4 clone37 (.A(net972),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(clknet_0_net470),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net40),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net1045),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(clknet_1_0__leaf_net289),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net55),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net919),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net940),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net295),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net785),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net954),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net1076),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net519),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net542),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net838),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net530),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net307),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net798),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net768),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net408),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net852),
    .X(net1164));
 sky130_fd_sc_hd__buf_12 fanout1 (.A(net969),
    .X(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap126_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c35_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A3 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_Y (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A4 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_B1_N (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_c48_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_X (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A0 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A2 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_S0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_Y (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A3 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_A1 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A1 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S1 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A1 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A3 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A3 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A3 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_c136_Y (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap104_A (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A3 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A1 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A1 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_Y (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_A2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_B1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_X (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SCD (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A3 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_D (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c139_X (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A2 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_A2 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A0 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A1 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c145_A2 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_X (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c144_A1 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer26_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_A1 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_X (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer20_A (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A3 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A2 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_A (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_A0 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_A2 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_X (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_A (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_B1 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_X (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap112_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A3 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_Y (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer4_A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_B1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A4 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_B1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c150_X (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_D (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S0 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_A (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A3 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_X (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A3 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A3 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_Y (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A4 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap74_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_Y (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCD (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_B1_N (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A4 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_A3 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A3 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c743_S0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c167_Y (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A3 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c168_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_SCD (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_D (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A3 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap97_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_Y (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_B1_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_A4 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A3 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A3 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_B1_N (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A3 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A3 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A4 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c184_Y (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_D (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCD (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A3 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A3 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A0 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A0 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A3 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A3 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_A3 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A3 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c180_A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A3 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c741_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_X (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A4 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_SCD (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_X (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_X (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A0 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A3 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCD (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_RESET_B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A0 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A1 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S1 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_X (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A3 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A3 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A4 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_Q_N (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A3 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_Q (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_B1_N (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_A3 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_A4 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_RESET_B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_B1_N (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap103_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A4 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_Y (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_Y (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c192_A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_S0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_c234_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap90_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_S1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_Y (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_A3 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_Q_N (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_Q (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net221_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A3 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_S0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_S1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A3 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_Y (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_X (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A3 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_Y (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A0 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_c269_Y (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap63_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_S0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_Y (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A3 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A0 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_c272_Y (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap56_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_A2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A3 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_c274_Y (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_A3 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_X (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c668_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_D (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_B1_N (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_Y (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A4 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_S0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_Y (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_S0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B1_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A3 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A2 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_S0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_D (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_RESET_B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A3 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SCD (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B1_N (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Q_N (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A0 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_Q (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_S1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c727_A0 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c703_A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A3 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_SCE (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_Y (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A3 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_Y (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_B1_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_D (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c300_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_X (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_c614_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_S0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A4 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_A0 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c296_Y (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_X (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_Y (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_D (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCD (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_SCE (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c369_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A4 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_B1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A3 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Q_N (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A3 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_A2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_Q (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c55_Y (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_SCD (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A3 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A3 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_B1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A4 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_Q (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold45_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_Q (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_S1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_Y (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c56_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_SCE (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A0 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_Q (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A3 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_Y (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A4 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A4 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net315_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_X (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_B1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A3 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_Y (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_S0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_Y (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_S0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_A3 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A0 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_RESET_B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_Y (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap57_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A0 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_Y (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A3 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A3 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_X (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_A1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_A4 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_X (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A0 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A0 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_A1 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_c404_Y (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_S0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_B1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_X (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_S0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A1 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SCE (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_RESET_B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_X (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A3 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A3 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SET_B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_X (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A3 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_D (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_X (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_B1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_A3 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SCD (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_X (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A3 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A3 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A2 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A3 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Q_N (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A3 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c415_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_A0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_Q (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_X (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_X (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_A0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A3 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c745_A3 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_S0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A2 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_D (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCE (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_X (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_SCE (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_SET_B (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_SCE (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_X (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_S0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A2 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_SCD (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c468_S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_B1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A4 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_A4 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A4 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_Q_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A3 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_A3 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_A3 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A3 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_Q (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCE (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A3 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_Q (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A2 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_X (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A3 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c426_Q (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A0 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A3 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c454_B1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_A3 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A3 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_A3 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A0 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A3 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_Q (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_X (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A3 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_A0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_X (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A2 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A3 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A0 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A0 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCE (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_X (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A0 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_SCD (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A0 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_Q (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c609_A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A3 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_S0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net456_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_X (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_A3 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_S0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_X (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net469_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_Y (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A3 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c355_A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_S0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c472_A3 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_B (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_X (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_A4 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_B (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_X (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_S0 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A0 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCE (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_B (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c532_X (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_Y (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A2 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A3 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_A4 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_Y (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A0 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_A2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_D (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c541_X (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c588_A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c542_Y (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_A3 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A0 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_RESET_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_RESET_B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c544_X (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_SCE (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_Q (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A0 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A0 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A4 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_X (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A3 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_A2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_X (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A3 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A3 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A0 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_A3 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCD (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_X (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_c98_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_Y (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A3 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_A0 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_A1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_X (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_c742_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A3 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_A4 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A3 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A4 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_X (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A2 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A2 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S0 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_X (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A3 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c705_A0 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_X (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_X (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_X (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_A0 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_S1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_SCD (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_D (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_X (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_X (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_S0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A3 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCE (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c39_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_Y (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_Y (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c516_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_X (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_S0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCD (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_X (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_A3 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_Y (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A3 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A0 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c744_A2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_X (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_A3 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_Y (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_B1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_A0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A0 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A3 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c675_X (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A3 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_X (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_A3 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SET_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_RESET_B (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_S0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_X (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_c719_S1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A2 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A2 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c690_A3 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_Q_N (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_A3 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c718_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A2 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_A2 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_Q (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_X (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_X (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_RESET_B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_X (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_D (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_X (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_D (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_X (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A4 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A4 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A3 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_S1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_S0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_c106_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_Q (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_Q (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c667_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c664_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c109_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold46_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_Q (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_S1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_Q (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_S0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_S0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_Q (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A3 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_S0 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_RESET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_Y (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_Q (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A3 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_S0 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_Q (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c553_B1_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_B1_N (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_c437_S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_Q (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A2 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S0 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c117_B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_S1 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B1_N (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_Q (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_B1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q_N (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_S1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_SCE (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_B1 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A4 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_Q (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c717_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_S1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A3 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_B1_N (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_Q (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_A3 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_Q (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A3 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c688_B1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_c659_S1 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_Q (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A2 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_Q (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A3 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S1 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_Q (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c766_S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c723_A2 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_A3 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_Q (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A3 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A2 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_Q (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_B1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c377_S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_S1 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_A3 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_Q (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c722_A3 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_S0 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_Q (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_S0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S1 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_Q (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A2 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_S0 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_Q (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A3 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_Q (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_A3 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c715_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S0 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_Q (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_S0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c503_S0 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_S1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_Q (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c502_S0 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A4 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q_N (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_S0 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_S1 (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_Q (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c525_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_Q (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_S1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A3 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_S0 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_s899_Q (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_Q (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c126_A4 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A3 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_Y (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net881_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_GCLK (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net882_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_GCLK (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_Q (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S0 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S1 (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_Q_N (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A3 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_S1 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_Q (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_A3 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_c363_S1 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_Q (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c724_A3 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c457_S1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c176_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q_N (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_S1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_Q (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_S1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c768_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c762_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c623_A3 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c476_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A3 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_Q (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_c590_S1 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_Q (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c733_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_S0 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_S1 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_A0 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_B1 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_X (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_A1 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A3 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_c625_S0 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_X (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c77_B (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c71_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c27_B (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A4 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A2 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_c123_A1 (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c769_A0 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c716_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c528_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_A2 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_A1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_S1 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_X (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A3 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c539_A1 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c33_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_B (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_A2 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_c28_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_S1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_B1 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_A3 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_c708_S0 (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_X (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A0 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_S1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A1 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c30_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_B (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A4 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A3 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_c202_B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_A0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S0 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c25_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A3 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_A2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c740_A2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c702_A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_S0 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_S1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c76_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c29_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_A1 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A3 (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c157_B (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_B1_N (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_A3 (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A4 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A2 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_S0 (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_A0 (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_B1_N (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_S0 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_c323_S1 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c90_Y (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S0 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A3 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap77_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c99_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_A3 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_Y (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_S1 (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_SCE (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A2 (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_X (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c635_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_A0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c655_A1 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c649_A3 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A2 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_X (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_Q (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A3 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c386_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_S0 (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_X (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_Y (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_S0 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_A3 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_A2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c629_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c493_A1 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A2 (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_X (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_S1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c262_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c259_A3 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c257_A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_X (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_X (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_RESET_B (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c709_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_A0 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_SCD (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_SCE (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_c589_A3 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_X (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c439_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A3 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_S0 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_A3 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_S0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_A0 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c494_A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A2 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_RESET_B (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_A3 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_S0 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A0 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_A3 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c756_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A2 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c765_A1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c760_S1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_SET_B (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_A2 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_SCD (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_A0 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A3 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A1 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c581_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_c628_A3 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_X (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c728_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_S0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A2 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c317_SET_B (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A3 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap56_X (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_S0 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A3 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c304_A2 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_S1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_c286_A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_S1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c293_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_B1_N (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c302_A4 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c292_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_B1 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c295_B1_N (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_c305_S0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_X (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_A4 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c435_B1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B1_N (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A4 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A2 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A3 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A3 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c487_A0 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_S1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_c350_A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer33_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A4 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_S1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A3 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_S1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_B1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap62_X (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c647_A0 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c513_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_A3 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap63_X (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_S0 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_A3 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_S1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c227_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A3 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_SCD (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_S0 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c207_S1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c361_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A0 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c195_A4 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_S1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_c243_A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A2 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_A3 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A0 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_X (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c384_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c383_A3 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c244_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_c235_A4 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_S0 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c225_A3 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c232_B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c165_B1_N (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c522_A0 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c249_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A3 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_S1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c86_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S0 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A3 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A4 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B1_N (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_S0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A0 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap74_X (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c646_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c492_S0 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c509_A1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_A3 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c621_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A3 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_S0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c228_A4 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_S0 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c105_B1_N (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_c100_B1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_X (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A3 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c63_S0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_A0 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap77_X (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_A0 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c504_A3 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c520_A1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_S1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_B1_N (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c61_B1_N (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c652_A0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_A3 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_S0 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_S1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A3 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c316_S0 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A3 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_SET_B (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A2 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_A1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_B1_N (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A4 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_S1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c707_S0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A0 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A3 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c84_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c258_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_S0 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A2 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A3 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_X (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c577_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_S1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_S1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_SCE (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c427_B1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A1 (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_SET_B (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_S1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c253_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A3 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_B1_N (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_S0 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_c191_A1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A0 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c488_A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c53_B1_N (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_B1_N (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c64_S1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_B1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c102_A1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B1_N (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_c60_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap89_X (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c653_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c624_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_B1 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_c91_B (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap90_X (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_S0 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c129_A4 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_c89_A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_X (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_S0 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_SCD (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c506_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_A3 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c194_A2 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_A1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_B1_N (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_X (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A4 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c389_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c368_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c263_S0 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c239_A3 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A2 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_c67_A (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_X (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c711_A1 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_S0 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A3 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_B (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_A1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_X (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c315_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_B1 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_S0 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_X (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c50_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_B (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap97_X (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c74_B (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_B (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A3 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_X (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c193_S1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c187_B1_N (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_B1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_S0 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c186_B1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_A3 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_A1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_B1_N (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap99_X (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c720_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c755_S0 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_c620_A2 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_X (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c412_B1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c406_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c408_S0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A3 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c757_A0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_S0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A1 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_S0 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap101_X (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_X (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_S0 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_B1_N (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_B1_N (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_A4 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap103_X (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c353_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c108_A1 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A2 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_X (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c691_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_A2 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge792_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_S0 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c569_A4 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_A3 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c563_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c560_S1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_SCD (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_B1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_X (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_S1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c747_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c730_A0 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_A2 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c591_A3 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_c575_A1 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_X (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c535_S0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c763_A3 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c761_S0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c749_S1 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A3 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c734_S1 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A2 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A0 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c407_B1_N (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_A4 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c446_A3 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c422_SCD (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A4 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SCE (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c411_B1_N (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_B1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_B1_N (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_X (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c698_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c684_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_B1_N (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_A4 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_A4 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A3 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_A2 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_c601_A1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_X (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c537_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c566_S1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S1 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_A3 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap112_X (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_A3 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_S0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_A1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_A1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_A1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A0 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_S1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap113_X (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c107_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c223_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c69_B (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_c40_B (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_A (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_S1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c93_B1_N (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c80_A4 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c70_A (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c256_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_A2 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c250_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A3 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A0 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c686_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c578_S0 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_B1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c451_B1_N (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_B1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_S1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c565_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c697_B1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_S1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_c699_B1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c559_B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c551_B1_N (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_SET_B (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c320_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_SCE (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_c306_S1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap120_X (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_S1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_A3 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c496_S0 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c291_A (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c421_B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c416_B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_c403_A (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_X (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c696_A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c459_A0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_S0 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_S1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c434_A4 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c432_A3 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c431_A1 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap123_X (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c118_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A2 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_c352_A4 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap124_X (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap123_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_B (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c51_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_c38_B1_N (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap125_X (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_A0 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_c31_A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap126_X (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c604_A2 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c485_S0 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c486_S1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_c92_B (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap127_X (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_A0 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c447_A2 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_B1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A4 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c584_S1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c313_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_B1_N (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_S0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_S0 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c526_A2 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_A1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_X (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c650_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c627_A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c603_A3 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c576_A3 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c533_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_S0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c182_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A2 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_c122_A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c657_A0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c517_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c507_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c73_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c379_S1 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c376_S0 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_SET_B (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_A4 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c198_A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_B1_N (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_A3 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_S0 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_c658_A2 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c97_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_RESET_B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c265_A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_A3 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c119_A1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c152_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c275_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_B1_N (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c94_A1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_S1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_SCE (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_S0 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_A3 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_B1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c764_A0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c693_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_A3 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c499_S0 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c471_A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c311_A4 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_B1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A2 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c26_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c190_A2 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_S0 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A0 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_A1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_c203_B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_A3 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_D (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c531_A1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c449_S0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A3 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_S0 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_A2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A3 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_S0 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c405_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c309_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c41_A4 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A0 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_A1 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_c143_B1_N (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_S0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c550_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c508_A0 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c260_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_S1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c169_A4 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_A1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c758_S0 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A0 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c420_A1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c521_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c428_A4 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c399_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c318_A3 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_A3 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c424_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c464_S0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S0 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c37_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c362_A3 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c34_B1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c78_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_A0 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A1 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c357_A3 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_SCE (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c208_B1_N (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B1_N (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c310_A3 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_S1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_B1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_B1_N (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c151_S0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_c149_S0 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c644_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c46_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_A2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_A1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_A3 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_B1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_X (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c158_B1_N (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c148_A2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c140_B1_N (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_B (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_B1_N (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c651_A1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c611_A0 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c600_A1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c582_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_A2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c400_B1_N (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c246_S0 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_B1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c179_A3 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_A1 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_S0 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c72_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c381_A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_S1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_A3 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c245_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c692_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c662_B (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A4 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c619_A0 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c62_A1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_A3 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c491_A2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c49_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_A4 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_A0 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_GATE_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_GATE (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge860_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s896_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s897_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s898_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c214_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_CLK_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c366_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge895_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GATE_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_SLEEP_B (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_GATE (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s905_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s918_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s945_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s946_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s944_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s956_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s960_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s961_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s940_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s955_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s957_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s958_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s959_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s933_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_GATE_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c423_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c556_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s949_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s950_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s951_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s952_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s953_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s954_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c548_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c669_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c681_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_GATE (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge862_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s947_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s948_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_S0 (.DIODE(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_A0 (.DIODE(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c714_S0 (.DIODE(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net567_X (.DIODE(clknet_1_1__leaf_net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_B1 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_S1 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_S0 (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net882_X (.DIODE(clknet_1_0__leaf_net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_c336_A3 (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c340_A3 (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_A3 (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c467_A0 (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A2 (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net313_X (.DIODE(clknet_1_1__leaf_net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_S1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A3 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_B1 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_S0 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c656_A2 (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net881_X (.DIODE(clknet_1_0__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_S1 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_S1 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_S0 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c605_S0 (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net881_X (.DIODE(clknet_1_1__leaf_net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_c319_D (.DIODE(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_A2 (.DIODE(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c456_A3 (.DIODE(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net289_X (.DIODE(clknet_1_1__leaf_net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_c205_A2 (.DIODE(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c222_A2 (.DIODE(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_A1 (.DIODE(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A4 (.DIODE(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net163_X (.DIODE(clknet_1_1__leaf_net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_c206_B1 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_S0 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c215_A1 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_S1 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_A3 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_S0 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_S1 (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net174_X (.DIODE(clknet_1_0__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c342_A4 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_A1 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_A2 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_A2 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c466_S0 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c490_A2 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_A2 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c630_A1 (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net174_X (.DIODE(clknet_1_1__leaf_net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_c345_SCD (.DIODE(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A2 (.DIODE(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_S0 (.DIODE(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net320_X (.DIODE(clknet_1_1__leaf_net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net177_A (.DIODE(clknet_0_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net177_A (.DIODE(clknet_0_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net177_X (.DIODE(clknet_0_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c209_A3 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A0 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A3 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A4 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_RESET_B (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c338_A4 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_S0 (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net177_X (.DIODE(clknet_1_0__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_A2 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_S0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c371_A0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_S0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c500_S0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A2 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S0 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c631_A1 (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net177_X (.DIODE(clknet_1_1__leaf_net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c210_A3 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c211_B1 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c212_A3 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_A3 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c216_A1 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c217_S0 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_A1 (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_SCD (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net178_X (.DIODE(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A1 (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_S1 (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A0 (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A1 (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_A3 (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net178_X (.DIODE(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_c221_A2 (.DIODE(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A1 (.DIODE(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c497_A1 (.DIODE(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net165_X (.DIODE(clknet_1_0__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c448_A3 (.DIODE(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c643_A0 (.DIODE(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c645_A3 (.DIODE(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c648_A3 (.DIODE(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net165_X (.DIODE(clknet_1_1__leaf_net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_A2 (.DIODE(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_c622_A0 (.DIODE(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net203_X (.DIODE(clknet_1_0__leaf_net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net161_A (.DIODE(clknet_0_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net161_A (.DIODE(clknet_0_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net161_X (.DIODE(clknet_0_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c322_A0 (.DIODE(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c450_A1 (.DIODE(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A2 (.DIODE(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net161_X (.DIODE(clknet_1_0__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_S0 (.DIODE(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A2 (.DIODE(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_S0 (.DIODE(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_c767_A0 (.DIODE(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net161_X (.DIODE(clknet_1_1__leaf_net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer3_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c397_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer2_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_X (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_X (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer14_A (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c665_A (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer13_A (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_X (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_A3 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A3 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_X (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_c737_A3 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_c752_A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer17_X (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer19_A (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_A0 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c616_S1 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c444_A2 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer18_X (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_c268_B1_N (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_B1_N (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c188_B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c199_A3 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_A4 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone30_X (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_c261_A0 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_A3 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c373_A3 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c236_B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone31_X (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_c701_S1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c251_S1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c618_A0 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_A1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_A3 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone32_X (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c173_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c254_S0 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c220_A1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone37_X (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c160_S0 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_S0 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c419_A3 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c418_A3 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c413_SCD (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone40_X (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_A0 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer42_X (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_X (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_c759_A2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c748_A1 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c695_A4 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone23_B1_N (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c54_B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c498_A2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c330_S0 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c185_A1 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_B1_N (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_B1_N (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net967));
 sky130_fd_sc_hd__mux4_1 clone1 (.A0(net1181),
    .A1(net1183),
    .A2(net1187),
    .A3(net1175),
    .S0(net1075),
    .S1(net1028),
    .X(net1166));
 sky130_fd_sc_hd__mux4_1 clone2 (.A0(net117),
    .A1(net1044),
    .A2(net1185),
    .A3(net1175),
    .S0(net1102),
    .S1(net1100),
    .X(net1167));
 sky130_fd_sc_hd__xnor2_1 clone3 (.A(net1075),
    .B(net105),
    .Y(net1168));
 sky130_fd_sc_hd__xnor2_1 clone4 (.A(net968),
    .B(net1075),
    .Y(net1169));
 sky130_fd_sc_hd__mux4_1 clone5 (.A0(net15),
    .A1(net9),
    .A2(net1056),
    .A3(net1052),
    .S0(net13),
    .S1(net1097),
    .X(net1170));
 sky130_fd_sc_hd__a31o_1 clone6 (.A1(net1092),
    .A2(net1088),
    .A3(net0),
    .B1(net1094),
    .X(net1171));
 sky130_fd_sc_hd__a21bo_1 clone7 (.A1(net108),
    .A2(net105),
    .B1_N(net1184),
    .X(net1172));
 sky130_fd_sc_hd__a31o_1 clone8 (.A1(net1092),
    .A2(net1088),
    .A3(net0),
    .B1(net1094),
    .X(net1173));
 sky130_fd_sc_hd__a21bo_1 clone9 (.A1(net1175),
    .A2(net1184),
    .B1_N(net1087),
    .X(net1174));
 sky130_fd_sc_hd__xnor2_1 clone10 (.A(net1075),
    .B(net105),
    .Y(net1175));
 sky130_fd_sc_hd__xnor2_1 clone11 (.A(net976),
    .B(net977),
    .Y(net1176));
 sky130_fd_sc_hd__a21bo_1 clone12 (.A1(net968),
    .A2(net1054),
    .B1_N(net1104),
    .X(net1177));
 sky130_fd_sc_hd__mux4_1 clone13 (.A0(net54),
    .A1(net56),
    .A2(net1031),
    .A3(net1046),
    .S0(net18),
    .S1(net979),
    .X(net1178));
 sky130_fd_sc_hd__mux4_1 clone14 (.A0(net118),
    .A1(net1183),
    .A2(net113),
    .A3(net106),
    .S0(net1075),
    .S1(net1028),
    .X(net1179));
 sky130_fd_sc_hd__a31o_1 clone15 (.A1(net120),
    .A2(net121),
    .A3(net1092),
    .B1(net1028),
    .X(net1180));
 sky130_fd_sc_hd__a41o_1 clone16 (.A1(net117),
    .A2(net1104),
    .A3(net103),
    .A4(net1039),
    .B1(net1042),
    .X(net1181));
 sky130_fd_sc_hd__a21bo_1 clone17 (.A1(net968),
    .A2(net1054),
    .B1_N(net1104),
    .X(net1182));
 sky130_fd_sc_hd__a31o_1 clone18 (.A1(net110),
    .A2(net113),
    .A3(net1044),
    .B1(net1063),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(net107),
    .X(net1184));
 sky130_fd_sc_hd__a41o_1 clone20 (.A1(net117),
    .A2(net1104),
    .A3(net103),
    .A4(net1039),
    .B1(net1042),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(net113),
    .X(net1186));
 sky130_fd_sc_hd__a21bo_1 clone24 (.A1(net1044),
    .A2(net106),
    .B1_N(net1097),
    .X(net1187));
 sky130_fd_sc_hd__clkbuf_1 clone25 (.A(net123),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(net969),
    .X(net1189));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
