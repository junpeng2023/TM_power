module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in25,
    in26,
    in27,
    in28,
    in29,
    in3,
    in30,
    in31,
    in32,
    in33,
    in34,
    in35,
    in36,
    in37,
    in38,
    in39,
    in4,
    in40,
    in41,
    in42,
    in43,
    in44,
    in45,
    in46,
    in47,
    in48,
    in49,
    in5,
    in50,
    in51,
    in52,
    in53,
    in54,
    in55,
    in56,
    in57,
    in58,
    in59,
    in6,
    in60,
    in61,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out25,
    out26,
    out27,
    out28,
    out29,
    out3,
    out30,
    out31,
    out32,
    out33,
    out34,
    out35,
    out36,
    out37,
    out38,
    out39,
    out4,
    out40,
    out41,
    out42,
    out43,
    out44,
    out45,
    out46,
    out47,
    out48,
    out49,
    out5,
    out50,
    out51,
    out52,
    out53,
    out54,
    out55,
    out56,
    out57,
    out58,
    out59,
    out6,
    out60,
    out61,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in25;
 input in26;
 input in27;
 input in28;
 input in29;
 input in3;
 input in30;
 input in31;
 input in32;
 input in33;
 input in34;
 input in35;
 input in36;
 input in37;
 input in38;
 input in39;
 input in4;
 input in40;
 input in41;
 input in42;
 input in43;
 input in44;
 input in45;
 input in46;
 input in47;
 input in48;
 input in49;
 input in5;
 input in50;
 input in51;
 input in52;
 input in53;
 input in54;
 input in55;
 input in56;
 input in57;
 input in58;
 input in59;
 input in6;
 input in60;
 input in61;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out25;
 output out26;
 output out27;
 output out28;
 output out29;
 output out3;
 output out30;
 output out31;
 output out32;
 output out33;
 output out34;
 output out35;
 output out36;
 output out37;
 output out38;
 output out39;
 output out4;
 output out40;
 output out41;
 output out42;
 output out43;
 output out44;
 output out45;
 output out46;
 output out47;
 output out48;
 output out49;
 output out5;
 output out50;
 output out51;
 output out52;
 output out53;
 output out54;
 output out55;
 output out56;
 output out57;
 output out58;
 output out59;
 output out6;
 output out60;
 output out61;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net679;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_net726;
 wire clknet_1_0__leaf_net726;
 wire clknet_1_1__leaf_net726;
 wire clknet_0_net808;
 wire clknet_1_0__leaf_net808;
 wire clknet_1_1__leaf_net808;
 wire clknet_0_net539;
 wire clknet_1_0__leaf_net539;
 wire clknet_1_1__leaf_net539;
 wire clknet_0_net553;
 wire clknet_1_0__leaf_net553;
 wire clknet_1_1__leaf_net553;
 wire clknet_0_net540;
 wire clknet_1_0__leaf_net540;
 wire clknet_1_1__leaf_net540;
 wire clknet_0_net725;
 wire clknet_1_0__leaf_net725;
 wire clknet_1_1__leaf_net725;
 wire clknet_0_net805;
 wire clknet_1_0__leaf_net805;
 wire clknet_1_1__leaf_net805;
 wire clknet_0_net424;
 wire clknet_1_0__leaf_net424;
 wire clknet_1_1__leaf_net424;
 wire clknet_0_net803;
 wire clknet_1_0__leaf_net803;
 wire clknet_1_1__leaf_net803;
 wire clknet_0_net422;
 wire clknet_1_0__leaf_net422;
 wire clknet_1_1__leaf_net422;
 wire clknet_0_net426;
 wire clknet_1_0__leaf_net426;
 wire clknet_1_1__leaf_net426;
 wire clknet_0_net813;
 wire clknet_1_0__leaf_net813;
 wire clknet_1_1__leaf_net813;
 wire clknet_0_net708;
 wire clknet_1_0__leaf_net708;
 wire clknet_1_1__leaf_net708;
 wire clknet_0_net306;
 wire clknet_1_0__leaf_net306;
 wire clknet_1_1__leaf_net306;
 wire clknet_0_net316;
 wire clknet_1_0__leaf_net316;
 wire clknet_1_1__leaf_net316;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net819;
 wire clknet_1_0__leaf_net819;
 wire clknet_1_1__leaf_net819;
 wire clknet_0_net198;
 wire clknet_1_0__leaf_net198;
 wire clknet_1_1__leaf_net198;
 wire clknet_0_net200;
 wire clknet_1_0__leaf_net200;
 wire clknet_1_1__leaf_net200;
 wire clknet_0_net199;
 wire clknet_1_0__leaf_net199;
 wire clknet_1_1__leaf_net199;
 wire clknet_0_net707;
 wire clknet_1_0__leaf_net707;
 wire clknet_1_1__leaf_net707;
 wire clknet_0_net660;
 wire clknet_1_0__leaf_net660;
 wire clknet_1_1__leaf_net660;
 wire clknet_0_net669;
 wire clknet_1_0__leaf_net669;
 wire clknet_1_1__leaf_net669;
 wire clknet_0_net661;
 wire clknet_1_0__leaf_net661;
 wire clknet_1_1__leaf_net661;
 wire clknet_0_net653;
 wire clknet_1_0__leaf_net653;
 wire clknet_1_1__leaf_net653;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net658;
 wire clknet_1_0__leaf_net658;
 wire clknet_1_1__leaf_net658;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net654;
 wire clknet_1_0__leaf_net654;
 wire clknet_1_1__leaf_net654;
 wire clknet_0_net656;
 wire clknet_1_0__leaf_net656;
 wire clknet_1_1__leaf_net656;
 wire clknet_0_net659;
 wire clknet_1_0__leaf_net659;
 wire clknet_1_1__leaf_net659;
 wire clknet_0_net652;
 wire clknet_1_0__leaf_net652;
 wire clknet_1_1__leaf_net652;
 wire clknet_0_net495;
 wire clknet_1_0__leaf_net495;
 wire clknet_1_1__leaf_net495;
 wire clknet_0_net493;
 wire clknet_1_0__leaf_net493;
 wire clknet_1_1__leaf_net493;
 wire clknet_0_net494;
 wire clknet_1_0__leaf_net494;
 wire clknet_1_1__leaf_net494;
 wire clknet_0_net292;
 wire clknet_1_0__leaf_net292;
 wire clknet_1_1__leaf_net292;
 wire clknet_0_net298;
 wire clknet_1_0__leaf_net298;
 wire clknet_1_1__leaf_net298;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net293;
 wire clknet_1_0__leaf_net293;
 wire clknet_1_1__leaf_net293;
 wire clknet_0_net294;
 wire clknet_1_0__leaf_net294;
 wire clknet_1_1__leaf_net294;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;

 sky130_fd_sc_hd__sdfxtp_1 c100 (.CLK(clknet_leaf_32_clk),
    .D(net867),
    .SCD(net929),
    .SCE(net36),
    .Q(net45));
 sky130_fd_sc_hd__sdfbbn_1 c101 (.CLK_N(clknet_leaf_32_clk),
    .D(net36),
    .RESET_B(net45),
    .SCD(net44),
    .SCE(net29),
    .SET_B(net35),
    .Q(net47),
    .Q_N(net46));
 sky130_fd_sc_hd__mux4_1 c102 (.A0(net37),
    .A1(net44),
    .A2(net45),
    .A3(net46),
    .S0(net27),
    .S1(net29),
    .X(net48));
 sky130_fd_sc_hd__sdfbbn_1 c103 (.CLK_N(clknet_leaf_32_clk),
    .D(net899),
    .RESET_B(net48),
    .SCD(net27),
    .SCE(net26),
    .SET_B(net35),
    .Q(net49));
 sky130_fd_sc_hd__a41o_1 c104 (.A1(net41),
    .A2(net49),
    .A3(net47),
    .A4(net43),
    .B1(net849),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 c105 (.A(net35),
    .X(net51));
 sky130_fd_sc_hd__buf_2 c106 (.A(net51),
    .X(net52));
 sky130_fd_sc_hd__xnor2_4 c107 (.A(net52),
    .B(net51),
    .Y(net53));
 sky130_fd_sc_hd__clkbuf_2 c108 (.A(net877),
    .X(net54));
 sky130_fd_sc_hd__xnor2_1 c109 (.A(net51),
    .B(net54),
    .Y(net55));
 sky130_fd_sc_hd__sdfxtp_1 c110 (.CLK(clknet_leaf_32_clk),
    .D(net51),
    .SCD(net54),
    .SCE(net53),
    .Q(net56));
 sky130_fd_sc_hd__a21bo_1 c111 (.A1(net952),
    .A2(net52),
    .B1_N(net54),
    .X(net57));
 sky130_fd_sc_hd__sdfxtp_1 c112 (.CLK(clknet_leaf_32_clk),
    .D(net52),
    .SCD(net54),
    .SCE(net53),
    .Q(net58));
 sky130_fd_sc_hd__clkbuf_2 c113 (.A(net686),
    .X(net59));
 sky130_fd_sc_hd__dfbbn_1 c114 (.CLK_N(clknet_leaf_31_clk),
    .D(net58),
    .RESET_B(net55),
    .SET_B(net53),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__dfbbn_1 c115 (.CLK_N(clknet_leaf_31_clk),
    .D(net55),
    .RESET_B(net53),
    .SET_B(net59),
    .Q(net63),
    .Q_N(net62));
 sky130_fd_sc_hd__a21bo_1 c116 (.A1(net56),
    .A2(net59),
    .B1_N(net51),
    .X(net814));
 sky130_fd_sc_hd__a21bo_1 c117 (.A1(net63),
    .A2(net59),
    .B1_N(net814),
    .X(net64));
 sky130_fd_sc_hd__dfbbp_1 c118 (.CLK(clknet_leaf_31_clk),
    .D(net57),
    .RESET_B(net64),
    .SET_B(net54),
    .Q(net66),
    .Q_N(net65));
 sky130_fd_sc_hd__a21bo_1 c119 (.A1(net59),
    .A2(net62),
    .B1_N(net54),
    .X(net67));
 sky130_fd_sc_hd__a21bo_1 c120 (.A1(net67),
    .A2(net66),
    .B1_N(net60),
    .X(net68));
 sky130_fd_sc_hd__sdfxbp_1 c121 (.CLK(clknet_leaf_31_clk),
    .D(net64),
    .SCD(net814),
    .SCE(net67),
    .Q(net70),
    .Q_N(net69));
 sky130_fd_sc_hd__mux4_1 c122 (.A0(net54),
    .A1(net67),
    .A2(net68),
    .A3(net65),
    .S0(net59),
    .S1(net51),
    .X(net71));
 sky130_fd_sc_hd__sdfxbp_1 c123 (.CLK(clknet_leaf_31_clk),
    .D(net68),
    .SCD(net71),
    .SCE(net67),
    .Q(net73),
    .Q_N(net72));
 sky130_fd_sc_hd__sdfxtp_1 c124 (.CLK(clknet_leaf_26_clk),
    .D(net71),
    .SCD(net61),
    .SCE(net910),
    .Q(net74));
 sky130_fd_sc_hd__mux4_1 c125 (.A0(net73),
    .A1(net70),
    .A2(net68),
    .A3(net74),
    .S0(net56),
    .S1(net52),
    .X(net75));
 sky130_fd_sc_hd__xnor2_4 c126 (.A(net745),
    .B(net760),
    .Y(net76));
 sky130_fd_sc_hd__xnor2_2 c127 (.A(net749),
    .B(net743),
    .Y(net77));
 sky130_fd_sc_hd__xnor2_1 c128 (.A(net76),
    .B(net750),
    .Y(net78));
 sky130_fd_sc_hd__a31o_1 c129 (.A1(net76),
    .A2(net78),
    .A3(net747),
    .B1(net77),
    .X(net79));
 sky130_fd_sc_hd__xnor2_1 c130 (.A(net76),
    .B(net748),
    .Y(net80));
 sky130_fd_sc_hd__sdfxtp_1 c131 (.CLK(clknet_leaf_7_clk),
    .D(net742),
    .SCD(net77),
    .SCE(net79),
    .Q(net81));
 sky130_fd_sc_hd__a21bo_1 c132 (.A1(net77),
    .A2(net781),
    .B1_N(net76),
    .X(net82));
 sky130_fd_sc_hd__sdfbbp_1 c133 (.CLK(clknet_leaf_7_clk),
    .D(net82),
    .RESET_B(net79),
    .SCD(net739),
    .SCE(net905),
    .SET_B(net76),
    .Q(net84),
    .Q_N(net83));
 sky130_fd_sc_hd__a21bo_1 c134 (.A1(net81),
    .A2(net679),
    .B1_N(net797),
    .X(net85));
 sky130_fd_sc_hd__xnor2_1 c135 (.A(net84),
    .B(net77),
    .Y(net86));
 sky130_fd_sc_hd__a21bo_1 c136 (.A1(net86),
    .A2(net85),
    .B1_N(net795),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 c137 (.A(net675),
    .X(net88));
 sky130_fd_sc_hd__a41o_1 c138 (.A1(net85),
    .A2(net77),
    .A3(net873),
    .A4(net86),
    .B1(net76),
    .X(net89));
 sky130_fd_sc_hd__sdfxtp_1 c139 (.CLK(clknet_leaf_5_clk),
    .D(net87),
    .SCD(net792),
    .SCE(net770),
    .Q(net90));
 sky130_fd_sc_hd__dfbbn_1 c140 (.CLK_N(clknet_leaf_5_clk),
    .D(net89),
    .RESET_B(net88),
    .SET_B(net79),
    .Q(net92),
    .Q_N(net91));
 sky130_fd_sc_hd__xnor2_1 c141 (.A(net90),
    .B(net91),
    .Y(net93));
 sky130_fd_sc_hd__dfbbn_1 c142 (.CLK_N(clknet_leaf_5_clk),
    .D(net79),
    .RESET_B(net93),
    .SET_B(net76),
    .Q(net94));
 sky130_fd_sc_hd__xnor2_1 c143 (.A(net92),
    .B(net94),
    .Y(net95));
 sky130_fd_sc_hd__buf_1 c144 (.A(net675),
    .X(net96));
 sky130_fd_sc_hd__a31o_1 c145 (.A1(net93),
    .A2(net95),
    .A3(net82),
    .B1(net81),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net97),
    .A1(net82),
    .A2(net740),
    .A3(net738),
    .S0(net93),
    .S1(net76),
    .X(net98));
 sky130_fd_sc_hd__a21bo_1 c147 (.A1(net763),
    .A2(net753),
    .B1_N(net757),
    .X(net99));
 sky130_fd_sc_hd__xnor2_1 c148 (.A(net99),
    .B(net933),
    .Y(net100));
 sky130_fd_sc_hd__a21bo_1 c149 (.A1(net764),
    .A2(net762),
    .B1_N(net772),
    .X(net101));
 sky130_fd_sc_hd__xnor2_2 c150 (.A(net99),
    .B(net751),
    .Y(net102));
 sky130_fd_sc_hd__xnor2_4 c151 (.A(net769),
    .B(net756),
    .Y(net103));
 sky130_fd_sc_hd__a21bo_1 c152 (.A1(net99),
    .A2(net103),
    .B1_N(net768),
    .X(net104));
 sky130_fd_sc_hd__a31o_1 c153 (.A1(net104),
    .A2(net758),
    .A3(net771),
    .B1(net100),
    .X(net105));
 sky130_fd_sc_hd__buf_1 c154 (.A(net838),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 c155 (.A0(net101),
    .A1(net102),
    .A2(net767),
    .A3(net105),
    .S0(net103),
    .S1(net106),
    .X(net107));
 sky130_fd_sc_hd__buf_1 c156 (.A(net671),
    .X(net108));
 sky130_fd_sc_hd__a21bo_1 c157 (.A1(net108),
    .A2(net106),
    .B1_N(net101),
    .X(net109));
 sky130_fd_sc_hd__sdfrbp_1 c158 (.CLK(clknet_leaf_4_clk),
    .D(net766),
    .RESET_B(net106),
    .SCD(net102),
    .SCE(net105),
    .Q(net111),
    .Q_N(net110));
 sky130_fd_sc_hd__xnor2_2 c159 (.A(net103),
    .B(net111),
    .Y(net112));
 sky130_fd_sc_hd__dfbbp_1 c160 (.CLK(clknet_leaf_0_clk),
    .D(net102),
    .RESET_B(net112),
    .SET_B(net105),
    .Q(net114),
    .Q_N(net113));
 sky130_fd_sc_hd__a21bo_1 c161 (.A1(net106),
    .A2(net108),
    .B1_N(net754),
    .X(net115));
 sky130_fd_sc_hd__a31o_1 c162 (.A1(net115),
    .A2(net110),
    .A3(net102),
    .B1(net112),
    .X(net116));
 sky130_fd_sc_hd__sdfxbp_1 c163 (.CLK(clknet_leaf_4_clk),
    .D(net100),
    .SCD(net116),
    .SCE(net112),
    .Q(net118),
    .Q_N(net117));
 sky130_fd_sc_hd__sdfrtn_1 c164 (.CLK_N(clknet_leaf_4_clk),
    .D(net111),
    .RESET_B(net116),
    .SCD(net112),
    .SCE(net117),
    .Q(net119));
 sky130_fd_sc_hd__a31o_1 c165 (.A1(net752),
    .A2(net843),
    .A3(net112),
    .B1(net119),
    .X(net120));
 sky130_fd_sc_hd__sdfrtp_1 c166 (.CLK(clknet_leaf_0_clk),
    .D(net108),
    .RESET_B(net844),
    .SCD(net116),
    .SCE(net103),
    .Q(net121));
 sky130_fd_sc_hd__mux4_1 c167 (.A0(net109),
    .A1(net114),
    .A2(net941),
    .A3(net120),
    .S0(net112),
    .S1(net103),
    .X(net122));
 sky130_fd_sc_hd__xnor2_4 c168 (.A(net0),
    .B(net774),
    .Y(net123));
 sky130_fd_sc_hd__xnor2_2 c169 (.A(net123),
    .B(net777),
    .Y(net124));
 sky130_fd_sc_hd__xnor2_1 c170 (.A(net123),
    .B(net776),
    .Y(net125));
 sky130_fd_sc_hd__dfstp_1 c171 (.CLK(clknet_leaf_35_clk),
    .D(net124),
    .SET_B(net125),
    .Q(net126));
 sky130_fd_sc_hd__sdfxbp_1 c172 (.CLK(clknet_leaf_35_clk),
    .D(net779),
    .SCD(net126),
    .SCE(net124),
    .Q(net128),
    .Q_N(net127));
 sky130_fd_sc_hd__xnor2_1 c173 (.A(net851),
    .B(net896),
    .Y(net129));
 sky130_fd_sc_hd__xnor2_2 c174 (.A(net123),
    .B(net851),
    .Y(net130));
 sky130_fd_sc_hd__xnor2_1 c175 (.A(net126),
    .B(net127),
    .Y(net131));
 sky130_fd_sc_hd__dfstp_1 c176 (.CLK(clknet_leaf_35_clk),
    .D(net896),
    .SET_B(net130),
    .Q(net132));
 sky130_fd_sc_hd__a31o_1 c177 (.A1(net786),
    .A2(net132),
    .A3(net126),
    .B1(net127),
    .X(net133));
 sky130_fd_sc_hd__a21bo_1 c178 (.A1(net129),
    .A2(net793),
    .B1_N(net131),
    .X(net134));
 sky130_fd_sc_hd__a21bo_1 c179 (.A1(net119),
    .A2(net129),
    .B1_N(net134),
    .X(net135));
 sky130_fd_sc_hd__sdfxtp_1 c180 (.CLK(clknet_leaf_35_clk),
    .D(net135),
    .SCD(net134),
    .SCE(net130),
    .Q(net136));
 sky130_fd_sc_hd__sdfxtp_1 c181 (.CLK(clknet_leaf_0_clk),
    .D(net887),
    .SCD(net135),
    .SCE(net131),
    .Q(net137));
 sky130_fd_sc_hd__sdfxtp_1 c182 (.CLK(clknet_leaf_35_clk),
    .D(net133),
    .SCD(net904),
    .SCE(net135),
    .Q(net138));
 sky130_fd_sc_hd__sdfrtp_1 c183 (.CLK(clknet_leaf_35_clk),
    .D(net125),
    .RESET_B(net852),
    .SCD(net138),
    .SCE(net904),
    .Q(net139));
 sky130_fd_sc_hd__a31o_1 c184 (.A1(net139),
    .A2(net133),
    .A3(net137),
    .B1(net138),
    .X(net140));
 sky130_fd_sc_hd__sdfrtp_1 c185 (.CLK(clknet_leaf_35_clk),
    .D(net130),
    .RESET_B(net135),
    .SCD(net140),
    .SCE(net138),
    .Q(net141));
 sky130_fd_sc_hd__a41o_1 c186 (.A1(net131),
    .A2(net138),
    .A3(net858),
    .A4(net137),
    .B1(net140),
    .X(net142));
 sky130_fd_sc_hd__sdfsbp_1 c187 (.CLK(clknet_leaf_35_clk),
    .D(net851),
    .SCD(net858),
    .SCE(net887),
    .SET_B(net859),
    .Q(net143));
 sky130_fd_sc_hd__sdfbbn_1 c188 (.CLK_N(clknet_leaf_35_clk),
    .D(net143),
    .RESET_B(net140),
    .SCD(net138),
    .SCE(net142),
    .SET_B(net124),
    .Q(net144));
 sky130_fd_sc_hd__buf_4 c189 (.A(net24),
    .X(net145));
 sky130_fd_sc_hd__buf_2 c190 (.A(net145),
    .X(net146));
 sky130_fd_sc_hd__xnor2_4 c191 (.A(net145),
    .B(net146),
    .Y(net147));
 sky130_fd_sc_hd__buf_1 c192 (.X(net681));
 sky130_fd_sc_hd__xnor2_1 c193 (.A(net146),
    .B(net145),
    .Y(net149));
 sky130_fd_sc_hd__clkbuf_1 c194 (.A(net680),
    .X(net150));
 sky130_fd_sc_hd__dfstp_2 c195 (.CLK(clknet_leaf_30_clk),
    .D(net150),
    .SET_B(net147),
    .Q(net151));
 sky130_fd_sc_hd__dlrbn_1 c196 (.D(net142),
    .GATE_N(clknet_leaf_1_clk),
    .RESET_B(net147),
    .Q(net153),
    .Q_N(net152));
 sky130_fd_sc_hd__a21bo_1 c197 (.A1(net148),
    .A2(net151),
    .B1_N(net150),
    .X(net154));
 sky130_fd_sc_hd__dfbbn_1 c198 (.CLK_N(clknet_leaf_1_clk),
    .D(net154),
    .RESET_B(net149),
    .SET_B(net151),
    .Q(net156),
    .Q_N(net155));
 sky130_fd_sc_hd__dlrbn_1 c199 (.D(net156),
    .GATE_N(clknet_leaf_30_clk),
    .RESET_B(net147),
    .Q(net158),
    .Q_N(net157));
 sky130_fd_sc_hd__xnor2_2 c200 (.A(net154),
    .B(net151),
    .Y(net159));
 sky130_fd_sc_hd__a21bo_1 c201 (.A1(net153),
    .A2(net159),
    .B1_N(net158),
    .X(net160));
 sky130_fd_sc_hd__a21bo_1 c202 (.A1(net158),
    .A2(net151),
    .B1_N(net148),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 c203 (.A0(net156),
    .A1(net158),
    .A2(net160),
    .A3(net147),
    .S0(net146),
    .S1(net145),
    .X(net162));
 sky130_fd_sc_hd__xnor2_1 c204 (.A(net151),
    .B(net159),
    .Y(net163));
 sky130_fd_sc_hd__mux4_1 c205 (.A0(net147),
    .A1(net163),
    .A2(net159),
    .A3(net155),
    .S0(net152),
    .S1(net157),
    .X(net164));
 sky130_fd_sc_hd__dfbbn_1 c206 (.CLK_N(clknet_leaf_1_clk),
    .D(net149),
    .RESET_B(net159),
    .SET_B(net939),
    .Q(net165));
 sky130_fd_sc_hd__dfbbp_1 c207 (.CLK(clknet_leaf_29_clk),
    .D(net146),
    .RESET_B(net163),
    .SET_B(net147),
    .Q(net167),
    .Q_N(net166));
 sky130_fd_sc_hd__mux4_1 c208 (.A0(net161),
    .A1(net165),
    .A2(net166),
    .A3(net157),
    .S0(net155),
    .S1(clknet_1_0__leaf_net707),
    .X(net168));
 sky130_fd_sc_hd__a21bo_1 c209 (.A1(net168),
    .A2(net706),
    .B1_N(clknet_1_1__leaf_net707),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 c210 (.A(net144),
    .X(net170));
 sky130_fd_sc_hd__xnor2_4 c211 (.A(net170),
    .B(net145),
    .Y(net171));
 sky130_fd_sc_hd__xnor2_1 c212 (.A(net170),
    .B(net171),
    .Y(net172));
 sky130_fd_sc_hd__xnor2_2 c213 (.A(net170),
    .B(net171),
    .Y(net173));
 sky130_fd_sc_hd__clkbuf_1 c214 (.A(net698),
    .X(net174));
 sky130_fd_sc_hd__xnor2_2 c215 (.A(net50),
    .B(net171),
    .Y(net175));
 sky130_fd_sc_hd__clkbuf_1 c216 (.A(net698),
    .X(net176));
 sky130_fd_sc_hd__sdfxbp_1 c217 (.CLK(clknet_leaf_30_clk),
    .D(net171),
    .SCD(net172),
    .SCE(net170),
    .Q(net178),
    .Q_N(net177));
 sky130_fd_sc_hd__dlrbp_1 c218 (.D(net178),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net173),
    .Q(net180),
    .Q_N(net179));
 sky130_fd_sc_hd__xnor2_1 c219 (.A(net176),
    .B(net177),
    .Y(net181));
 sky130_fd_sc_hd__dlrbp_1 c220 (.D(net180),
    .GATE(clknet_leaf_30_clk),
    .RESET_B(net172),
    .Q(net183),
    .Q_N(net182));
 sky130_fd_sc_hd__a21bo_2 c221 (.A1(net181),
    .A2(net855),
    .B1_N(net170),
    .X(net184));
 sky130_fd_sc_hd__a21bo_1 c222 (.A1(net174),
    .A2(net180),
    .B1_N(net184),
    .X(net185));
 sky130_fd_sc_hd__xnor2_2 c223 (.A(net184),
    .B(net906),
    .Y(net186));
 sky130_fd_sc_hd__dlrtn_1 c224 (.D(net185),
    .GATE_N(clknet_leaf_31_clk),
    .RESET_B(net186),
    .Q(net187));
 sky130_fd_sc_hd__sdfsbp_1 c225 (.CLK(clknet_leaf_31_clk),
    .D(net187),
    .SCD(net173),
    .SCE(net170),
    .SET_B(net171),
    .Q(net189),
    .Q_N(net188));
 sky130_fd_sc_hd__sdfstp_1 c226 (.CLK(clknet_leaf_29_clk),
    .D(net173),
    .SCD(net171),
    .SCE(net897),
    .SET_B(net856),
    .Q(net190));
 sky130_fd_sc_hd__dlrtn_1 c227 (.D(net913),
    .GATE_N(clknet_leaf_26_clk),
    .RESET_B(net186),
    .Q(net191));
 sky130_fd_sc_hd__sdfxbp_1 c228 (.CLK(clknet_leaf_29_clk),
    .D(net881),
    .SCD(net184),
    .SCE(net185),
    .Q(net192));
 sky130_fd_sc_hd__a41o_1 c229 (.A1(net183),
    .A2(net192),
    .A3(net188),
    .A4(net184),
    .B1(net171),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 c230 (.A0(net191),
    .A1(net193),
    .A2(net189),
    .A3(net184),
    .S0(net171),
    .S1(net173),
    .X(net194));
 sky130_fd_sc_hd__buf_4 c231 (.X(net195));
 sky130_fd_sc_hd__xnor2_1 c232 (.A(net827),
    .B(clknet_1_0__leaf_net708),
    .Y(net196));
 sky130_fd_sc_hd__xnor2_1 c233 (.A(net74),
    .B(net826),
    .Y(net197));
 sky130_fd_sc_hd__xnor2_1 c234 (.A(clknet_1_0__leaf_net196),
    .B(net827),
    .Y(net198));
 sky130_fd_sc_hd__a21bo_1 c235 (.A1(clknet_1_0__leaf_net198),
    .A2(net197),
    .B1_N(net826),
    .X(net199));
 sky130_fd_sc_hd__xnor2_1 c236 (.A(net826),
    .B(clknet_1_1__leaf_net198),
    .Y(net200));
 sky130_fd_sc_hd__clkbuf_1 c237 (.A(net678),
    .X(net201));
 sky130_fd_sc_hd__a21bo_1 c238 (.A1(net826),
    .A2(net197),
    .B1_N(net69),
    .X(net804));
 sky130_fd_sc_hd__mux4_1 c239 (.A0(net197),
    .A1(net804),
    .A2(clknet_1_1__leaf_net199),
    .A3(net826),
    .S0(clknet_1_0__leaf_net200),
    .S1(net69),
    .X(net202));
 sky130_fd_sc_hd__xnor2_4 c240 (.A(net827),
    .B(net709),
    .Y(net203));
 sky130_fd_sc_hd__mux4_1 c241 (.A0(clknet_1_0__leaf_net199),
    .A1(net804),
    .A2(net197),
    .A3(clknet_1_0__leaf_net200),
    .S0(net826),
    .S1(clknet_1_0__leaf_net198),
    .X(net204));
 sky130_fd_sc_hd__a41o_1 c242 (.A1(net201),
    .A2(net74),
    .A3(net826),
    .A4(net69),
    .B1(net710),
    .X(net205));
 sky130_fd_sc_hd__xnor2_4 c243 (.A(net70),
    .B(net203),
    .Y(net206));
 sky130_fd_sc_hd__a21bo_1 c244 (.A1(net206),
    .A2(net826),
    .B1_N(net711),
    .X(net207));
 sky130_fd_sc_hd__sdfxtp_1 c245 (.CLK(clknet_leaf_25_clk),
    .D(net207),
    .SCD(net205),
    .SCE(net827),
    .Q(net208));
 sky130_fd_sc_hd__sdfbbn_1 c246 (.CLK_N(clknet_leaf_26_clk),
    .D(net903),
    .RESET_B(net864),
    .SCD(net206),
    .SCE(net53),
    .SET_B(net175),
    .Q(net210),
    .Q_N(net209));
 sky130_fd_sc_hd__sdfxtp_1 c247 (.CLK(clknet_leaf_25_clk),
    .D(clknet_1_1__leaf_net200),
    .SCD(net891),
    .SCE(net826),
    .Q(net211));
 sky130_fd_sc_hd__mux4_2 c248 (.A0(net206),
    .A1(clknet_1_1__leaf_net196),
    .A2(net209),
    .A3(net208),
    .S0(net804),
    .S1(net827),
    .X(net819));
 sky130_fd_sc_hd__mux4_1 c249 (.A0(net210),
    .A1(net208),
    .A2(clknet_1_1__leaf_net199),
    .A3(net205),
    .S0(net70),
    .S1(net827),
    .X(net212));
 sky130_fd_sc_hd__sdfbbp_1 c250 (.CLK(clknet_leaf_25_clk),
    .D(net186),
    .RESET_B(net205),
    .SCD(net890),
    .SCE(clknet_1_1__leaf_net819),
    .SET_B(net845),
    .Q(net820),
    .Q_N(net213));
 sky130_fd_sc_hd__mux4_1 c251 (.A0(net205),
    .A1(net211),
    .A2(net213),
    .A3(net206),
    .S0(net826),
    .S1(clknet_1_1__leaf_net200),
    .X(net214));
 sky130_fd_sc_hd__dlymetal6s2s_1 c252 (.A(net96),
    .X(net215));
 sky130_fd_sc_hd__xnor2_2 c253 (.A(net215),
    .B(net746),
    .Y(net216));
 sky130_fd_sc_hd__a21bo_2 c254 (.A1(net216),
    .A2(net744),
    .B1_N(net215),
    .X(net217));
 sky130_fd_sc_hd__buf_1 c255 (.X(net218));
 sky130_fd_sc_hd__clkbuf_1 c256 (.A(net673),
    .X(net219));
 sky130_fd_sc_hd__dlrtn_2 c257 (.D(net216),
    .GATE_N(clknet_leaf_7_clk),
    .RESET_B(net217),
    .Q(net220));
 sky130_fd_sc_hd__dlrtp_1 c258 (.D(net217),
    .GATE(clknet_leaf_7_clk),
    .RESET_B(net216),
    .Q(net221));
 sky130_fd_sc_hd__a21bo_1 c259 (.A1(net796),
    .A2(net216),
    .B1_N(net220),
    .X(net222));
 sky130_fd_sc_hd__sdfxtp_1 c260 (.CLK(clknet_leaf_7_clk),
    .D(net78),
    .SCD(net222),
    .SCE(net220),
    .Q(net223));
 sky130_fd_sc_hd__dfbbn_1 c261 (.CLK_N(clknet_leaf_7_clk),
    .D(net215),
    .RESET_B(net901),
    .SET_B(net217),
    .Q(net224));
 sky130_fd_sc_hd__xnor2_1 c262 (.A(net224),
    .B(net223),
    .Y(net225));
 sky130_fd_sc_hd__dfbbn_1 c263 (.CLK_N(clknet_leaf_7_clk),
    .D(net217),
    .RESET_B(net901),
    .SET_B(net223),
    .Q(net227),
    .Q_N(net226));
 sky130_fd_sc_hd__a31o_1 c264 (.A1(net221),
    .A2(net227),
    .A3(net225),
    .B1(net220),
    .X(net228));
 sky130_fd_sc_hd__sdfstp_1 c265 (.CLK(clknet_leaf_7_clk),
    .D(net909),
    .SCD(net226),
    .SCE(net225),
    .SET_B(net217),
    .Q(net229));
 sky130_fd_sc_hd__a21bo_1 c266 (.A1(net219),
    .A2(net220),
    .B1_N(net218),
    .X(net230));
 sky130_fd_sc_hd__a21bo_1 c267 (.A1(net229),
    .A2(net218),
    .B1_N(net230),
    .X(net231));
 sky130_fd_sc_hd__mux4_1 c268 (.A0(net218),
    .A1(net225),
    .A2(net229),
    .A3(net231),
    .S0(net217),
    .S1(net220),
    .X(net232));
 sky130_fd_sc_hd__a21bo_1 c269 (.A1(net230),
    .A2(net229),
    .B1_N(net714),
    .X(net233));
 sky130_fd_sc_hd__a21bo_1 c270 (.A1(net227),
    .A2(net230),
    .B1_N(net233),
    .X(net234));
 sky130_fd_sc_hd__mux4_1 c271 (.A0(net220),
    .A1(net229),
    .A2(net233),
    .A3(net226),
    .S0(net231),
    .S1(net217),
    .X(net235));
 sky130_fd_sc_hd__mux4_1 c272 (.A0(net234),
    .A1(net233),
    .A2(net230),
    .A3(net220),
    .S0(net231),
    .S1(net715),
    .X(net236));
 sky130_fd_sc_hd__buf_4 c273 (.A(in32),
    .X(net237));
 sky130_fd_sc_hd__xnor2_4 c274 (.A(net237),
    .B(net716),
    .Y(net238));
 sky130_fd_sc_hd__xnor2_1 c275 (.A(net237),
    .B(net238),
    .Y(net239));
 sky130_fd_sc_hd__clkbuf_1 c276 (.X(net240));
 sky130_fd_sc_hd__buf_1 c277 (.A(net691),
    .X(net241));
 sky130_fd_sc_hd__a21bo_1 c278 (.A1(net241),
    .A2(net238),
    .B1_N(net237),
    .X(net242));
 sky130_fd_sc_hd__xnor2_1 c279 (.A(net241),
    .B(net755),
    .Y(net243));
 sky130_fd_sc_hd__a21bo_1 c280 (.A1(net243),
    .A2(net238),
    .B1_N(net237),
    .X(net244));
 sky130_fd_sc_hd__dfbbp_1 c281 (.CLK(clknet_leaf_4_clk),
    .D(net857),
    .RESET_B(net239),
    .SET_B(net237),
    .Q(net246),
    .Q_N(net245));
 sky130_fd_sc_hd__sdfxbp_1 c282 (.CLK(clknet_leaf_3_clk),
    .D(net242),
    .SCD(net246),
    .SCE(net918),
    .Q(net248),
    .Q_N(net247));
 sky130_fd_sc_hd__a21bo_1 c283 (.A1(net247),
    .A2(net246),
    .B1_N(net704),
    .X(net249));
 sky130_fd_sc_hd__a21bo_1 c284 (.A1(net238),
    .A2(net243),
    .B1_N(net249),
    .X(net250));
 sky130_fd_sc_hd__sdfxbp_1 c285 (.CLK(clknet_leaf_3_clk),
    .D(net244),
    .SCD(net246),
    .SCE(net249),
    .Q(net252),
    .Q_N(net251));
 sky130_fd_sc_hd__sdfxtp_1 c286 (.CLK(clknet_leaf_5_clk),
    .D(net239),
    .SCD(net244),
    .SCE(net246),
    .Q(net253));
 sky130_fd_sc_hd__sdfxtp_1 c287 (.CLK(clknet_leaf_5_clk),
    .D(net868),
    .SCD(net242),
    .SCE(net249),
    .Q(net254));
 sky130_fd_sc_hd__mux4_1 c288 (.A0(net233),
    .A1(net250),
    .A2(net254),
    .A3(net238),
    .S0(net245),
    .S1(net237),
    .X(net255));
 sky130_fd_sc_hd__a21bo_1 c289 (.A1(net249),
    .A2(net253),
    .B1_N(net761),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 c290 (.A0(net250),
    .A1(net958),
    .A2(net244),
    .A3(net238),
    .S0(net237),
    .S1(net256),
    .X(net257));
 sky130_fd_sc_hd__a21bo_1 c291 (.A1(net256),
    .A2(net237),
    .B1_N(net718),
    .X(net258));
 sky130_fd_sc_hd__sdfxtp_1 c292 (.CLK(clknet_leaf_6_clk),
    .D(net258),
    .SCD(net256),
    .SCE(net249),
    .Q(net259));
 sky130_fd_sc_hd__dfbbn_1 c293 (.CLK_N(clknet_leaf_6_clk),
    .D(net259),
    .RESET_B(net258),
    .SET_B(net719),
    .Q(net260));
 sky130_fd_sc_hd__xnor2_4 c294 (.A(net828),
    .B(net717),
    .Y(net261));
 sky130_fd_sc_hd__xnor2_4 c295 (.A(net261),
    .B(net245),
    .Y(net262));
 sky130_fd_sc_hd__xnor2_1 c296 (.A(net261),
    .B(net262),
    .Y(net263));
 sky130_fd_sc_hd__clkbuf_2 c297 (.A(net942),
    .X(net815));
 sky130_fd_sc_hd__xnor2_1 c298 (.A(net953),
    .B(net261),
    .Y(net264));
 sky130_fd_sc_hd__xnor2_2 c299 (.A(net815),
    .B(net262),
    .Y(net265));
 sky130_fd_sc_hd__buf_1 c300 (.A(net672),
    .X(net266));
 sky130_fd_sc_hd__dlrtp_1 c301 (.D(net265),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net266),
    .Q(net267));
 sky130_fd_sc_hd__dlrtp_1 c302 (.D(net264),
    .GATE(clknet_leaf_2_clk),
    .RESET_B(net265),
    .Q(net268));
 sky130_fd_sc_hd__edfxbp_1 c303 (.CLK(clknet_leaf_2_clk),
    .D(net263),
    .DE(net922),
    .Q(net270),
    .Q_N(net269));
 sky130_fd_sc_hd__a21bo_1 c304 (.A1(net268),
    .A2(net266),
    .B1_N(net267),
    .X(net271));
 sky130_fd_sc_hd__xnor2_2 c305 (.A(net267),
    .B(net853),
    .Y(net272));
 sky130_fd_sc_hd__a41o_1 c306 (.A1(net272),
    .A2(net270),
    .A3(net268),
    .A4(net266),
    .B1(net828),
    .X(net273));
 sky130_fd_sc_hd__dfbbn_1 c307 (.CLK_N(clknet_leaf_2_clk),
    .D(net266),
    .RESET_B(net268),
    .SET_B(net265),
    .Q(net275),
    .Q_N(net274));
 sky130_fd_sc_hd__a21bo_1 c308 (.A1(net273),
    .A2(net271),
    .B1_N(net269),
    .X(net276));
 sky130_fd_sc_hd__a21bo_1 c309 (.A1(net262),
    .A2(net274),
    .B1_N(net269),
    .X(net277));
 sky130_fd_sc_hd__a21bo_1 c310 (.A1(net275),
    .A2(net271),
    .B1_N(net267),
    .X(net278));
 sky130_fd_sc_hd__dfbbp_1 c311 (.CLK(clknet_leaf_2_clk),
    .D(net278),
    .RESET_B(net277),
    .SET_B(net854),
    .Q(net280),
    .Q_N(net279));
 sky130_fd_sc_hd__mux4_1 c312 (.A0(net267),
    .A1(net278),
    .A2(net272),
    .A3(net279),
    .S0(net273),
    .S1(net262),
    .X(net281));
 sky130_fd_sc_hd__sdfxbp_1 c313 (.CLK(clknet_leaf_2_clk),
    .D(net281),
    .SCD(net276),
    .SCE(net280),
    .Q(net283),
    .Q_N(net282));
 sky130_fd_sc_hd__sdfbbn_1 c314 (.CLK_N(clknet_leaf_2_clk),
    .D(net280),
    .RESET_B(net281),
    .SCD(net265),
    .SCE(net272),
    .SET_B(net261),
    .Q(net284));
 sky130_fd_sc_hd__clkbuf_2 c315 (.A(net283),
    .X(net285));
 sky130_fd_sc_hd__xnor2_1 c316 (.A(net283),
    .B(net285),
    .Y(net286));
 sky130_fd_sc_hd__edfxtp_1 c317 (.CLK(clknet_leaf_2_clk),
    .D(net277),
    .DE(net285),
    .Q(net287));
 sky130_fd_sc_hd__xnor2_1 c318 (.A(net270),
    .B(net287),
    .Y(net288));
 sky130_fd_sc_hd__xnor2_1 c319 (.A(net286),
    .B(net285),
    .Y(net289));
 sky130_fd_sc_hd__xnor2_1 c320 (.A(net285),
    .B(net287),
    .Y(net290));
 sky130_fd_sc_hd__xnor2_1 c321 (.A(net284),
    .B(net290),
    .Y(net291));
 sky130_fd_sc_hd__sdlclkp_1 c322 (.CLK(clknet_leaf_29_clk),
    .GATE(net145),
    .SCE(net291),
    .GCLK(net292));
 sky130_fd_sc_hd__xnor2_1 c323 (.A(net288),
    .B(clknet_1_1__leaf_net292),
    .Y(net293));
 sky130_fd_sc_hd__xnor2_1 c324 (.A(net287),
    .B(clknet_1_0__leaf_net293),
    .Y(net294));
 sky130_fd_sc_hd__sdfxbp_1 c325 (.CLK(clknet_leaf_29_clk),
    .D(net290),
    .SCD(clknet_1_0__leaf_net293),
    .SCE(clknet_1_1__leaf_net294),
    .Q(net296),
    .Q_N(net295));
 sky130_fd_sc_hd__sdfxtp_2 c326 (.CLK(clknet_leaf_29_clk),
    .D(clknet_1_0__leaf_net292),
    .SCD(net291),
    .SCE(clknet_1_0__leaf_net294),
    .Q(net297));
 sky130_fd_sc_hd__a21bo_1 c327 (.A1(net261),
    .A2(clknet_1_0__leaf_net292),
    .B1_N(net297),
    .X(net298));
 sky130_fd_sc_hd__sdlclkp_2 c328 (.CLK(clknet_leaf_29_clk),
    .GATE(clknet_1_0__leaf_net294),
    .SCE(net842),
    .GCLK(net299));
 sky130_fd_sc_hd__sdfxtp_2 c329 (.CLK(clknet_leaf_29_clk),
    .D(net160),
    .SCD(net842),
    .SCE(clknet_1_0__leaf_net298),
    .Q(net300));
 sky130_fd_sc_hd__sdfstp_1 c330 (.CLK(clknet_leaf_29_clk),
    .D(net291),
    .SCD(net961),
    .SCE(clknet_1_0__leaf_net298),
    .SET_B(net842),
    .Q(net818));
 sky130_fd_sc_hd__a31o_1 c331 (.A1(clknet_1_1__leaf_net298),
    .A2(net296),
    .A3(net297),
    .B1(net300),
    .X(net301));
 sky130_fd_sc_hd__sedfxbp_1 c332 (.CLK(clknet_leaf_29_clk),
    .D(net289),
    .DE(net299),
    .SCD(net923),
    .SCE(clknet_1_1__leaf_net301),
    .Q(net302));
 sky130_fd_sc_hd__sedfxbp_1 c333 (.CLK(clknet_leaf_28_clk),
    .D(net302),
    .DE(clknet_1_0__leaf_net301),
    .SCD(net961),
    .SCE(net818),
    .Q(net304),
    .Q_N(net303));
 sky130_fd_sc_hd__a31o_1 c334 (.A1(net167),
    .A2(net295),
    .A3(net300),
    .B1(net303),
    .X(net821));
 sky130_fd_sc_hd__xnor2_1 c335 (.A(clknet_1_1__leaf_net293),
    .B(net304),
    .Y(net305));
 sky130_fd_sc_hd__xnor2_2 c336 (.A(net296),
    .B(clknet_1_1__leaf_net708),
    .Y(net306));
 sky130_fd_sc_hd__buf_1 c337 (.A(clknet_1_0__leaf_net306),
    .X(net307));
 sky130_fd_sc_hd__xnor2_1 c338 (.A(clknet_1_1__leaf_net306),
    .B(clknet_1_1__leaf_net307),
    .Y(net308));
 sky130_fd_sc_hd__buf_2 c339 (.A(net683),
    .X(net309));
 sky130_fd_sc_hd__buf_1 c340 (.A(net682),
    .X(net310));
 sky130_fd_sc_hd__xnor2_1 c341 (.A(net309),
    .B(clknet_1_1__leaf_net307),
    .Y(net311));
 sky130_fd_sc_hd__xnor2_1 c342 (.A(clknet_1_0__leaf_net307),
    .B(net309),
    .Y(net312));
 sky130_fd_sc_hd__xnor2_2 c343 (.A(net842),
    .B(net309),
    .Y(net313));
 sky130_fd_sc_hd__sdlclkp_4 c344 (.CLK(clknet_leaf_28_clk),
    .GATE(net310),
    .SCE(net312),
    .GCLK(net314));
 sky130_fd_sc_hd__xnor2_2 c345 (.A(net313),
    .B(net309),
    .Y(net315));
 sky130_fd_sc_hd__a21bo_1 c346 (.A1(net314),
    .A2(clknet_1_0__leaf_net306),
    .B1_N(net309),
    .X(net316));
 sky130_fd_sc_hd__sdfxtp_1 c347 (.CLK(clknet_leaf_27_clk),
    .D(net311),
    .SCD(clknet_1_0__leaf_net316),
    .SCE(clknet_1_0__leaf_net306),
    .Q(net317));
 sky130_fd_sc_hd__xnor2_2 c348 (.A(net315),
    .B(net313),
    .Y(net318));
 sky130_fd_sc_hd__dfrbp_1 c349 (.CLK(clknet_leaf_27_clk),
    .D(clknet_1_0__leaf_net316),
    .RESET_B(net318),
    .Q(net319));
 sky130_fd_sc_hd__a21bo_1 c350 (.A1(net319),
    .A2(net317),
    .B1_N(clknet_1_1__leaf_net307),
    .X(net320));
 sky130_fd_sc_hd__dfbbn_1 c351 (.CLK_N(clknet_leaf_28_clk),
    .D(net318),
    .RESET_B(clknet_1_1__leaf_net306),
    .SET_B(clknet_1_1__leaf_net316),
    .Q(net322),
    .Q_N(net321));
 sky130_fd_sc_hd__dfbbn_1 c352 (.CLK_N(clknet_leaf_28_clk),
    .D(net308),
    .RESET_B(net317),
    .SET_B(net886),
    .Q(net324),
    .Q_N(net323));
 sky130_fd_sc_hd__sedfxtp_1 c353 (.CLK(clknet_leaf_27_clk),
    .D(net324),
    .DE(net320),
    .SCD(net318),
    .SCE(net310),
    .Q(net325));
 sky130_fd_sc_hd__a21bo_1 c354 (.A1(net322),
    .A2(net309),
    .B1_N(clknet_1_1__leaf_net306),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 c355 (.A0(net326),
    .A1(net315),
    .A2(net325),
    .A3(clknet_1_1__leaf_net316),
    .S0(net318),
    .S1(net321),
    .X(net327));
 sky130_fd_sc_hd__a21bo_1 c356 (.A1(net325),
    .A2(net323),
    .B1_N(net720),
    .X(net816));
 sky130_fd_sc_hd__xnor2_1 c377 (.A(net804),
    .B(net713),
    .Y(net817));
 sky130_fd_sc_hd__clkbuf_8 c378 (.A(net825),
    .X(net328));
 sky130_fd_sc_hd__xnor2_1 c379 (.A(net328),
    .B(net825),
    .Y(net329));
 sky130_fd_sc_hd__xnor2_1 c380 (.A(net228),
    .B(net328),
    .Y(net330));
 sky130_fd_sc_hd__clkbuf_1 c381 (.A(net694),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 c382 (.A(net954),
    .X(net332));
 sky130_fd_sc_hd__xnor2_1 c383 (.A(net331),
    .B(net332),
    .Y(net333));
 sky130_fd_sc_hd__xnor2_4 c384 (.A(net328),
    .B(net332),
    .Y(net334));
 sky130_fd_sc_hd__xnor2_2 c385 (.A(net334),
    .B(net328),
    .Y(net335));
 sky130_fd_sc_hd__dfrbp_1 c386 (.CLK(clknet_leaf_8_clk),
    .D(net334),
    .RESET_B(net335),
    .Q(net337),
    .Q_N(net336));
 sky130_fd_sc_hd__sedfxtp_4 c387 (.CLK(clknet_leaf_8_clk),
    .D(net332),
    .DE(net336),
    .SCD(net335),
    .SCE(net334),
    .Q(net338));
 sky130_fd_sc_hd__dfrtn_1 c388 (.CLK_N(clknet_leaf_9_clk),
    .D(net335),
    .RESET_B(net338),
    .Q(net339));
 sky130_fd_sc_hd__dfbbp_1 c389 (.CLK(clknet_leaf_8_clk),
    .D(net329),
    .RESET_B(net339),
    .SET_B(net335),
    .Q(net341),
    .Q_N(net340));
 sky130_fd_sc_hd__sdfxbp_2 c390 (.CLK(clknet_leaf_9_clk),
    .D(net339),
    .SCD(net335),
    .SCE(net338),
    .Q(net343),
    .Q_N(net342));
 sky130_fd_sc_hd__xnor2_1 c391 (.A(net337),
    .B(net338),
    .Y(net344));
 sky130_fd_sc_hd__a41o_1 c392 (.A1(net341),
    .A2(net343),
    .A3(net338),
    .A4(net334),
    .B1(net332),
    .X(net345));
 sky130_fd_sc_hd__sdfbbn_1 c393 (.CLK_N(clknet_leaf_8_clk),
    .D(net333),
    .RESET_B(net343),
    .SCD(net338),
    .SCE(net335),
    .SET_B(net332),
    .Q(net346));
 sky130_fd_sc_hd__a41o_1 c394 (.A1(net231),
    .A2(net344),
    .A3(net339),
    .A4(net343),
    .B1(net338),
    .X(net347));
 sky130_fd_sc_hd__sdfbbp_1 c395 (.CLK(clknet_leaf_9_clk),
    .D(net96),
    .RESET_B(net347),
    .SCD(net328),
    .SCE(net342),
    .SET_B(net332),
    .Q(net349),
    .Q_N(net348));
 sky130_fd_sc_hd__xnor2_1 c396 (.A(net349),
    .B(net340),
    .Y(net350));
 sky130_fd_sc_hd__xnor2_1 c397 (.A(net350),
    .B(net349),
    .Y(net351));
 sky130_fd_sc_hd__mux4_1 c398 (.A0(net346),
    .A1(net351),
    .A2(net350),
    .A3(net348),
    .S0(net342),
    .S1(net338),
    .X(net352));
 sky130_fd_sc_hd__xnor2_4 c399 (.A(net252),
    .B(net343),
    .Y(net353));
 sky130_fd_sc_hd__xnor2_2 c400 (.A(net260),
    .B(net353),
    .Y(net354));
 sky130_fd_sc_hd__xnor2_1 c401 (.A(net353),
    .B(net823),
    .Y(net355));
 sky130_fd_sc_hd__clkbuf_2 c402 (.A(net831),
    .X(net356));
 sky130_fd_sc_hd__xnor2_1 c403 (.A(net246),
    .B(net356),
    .Y(net357));
 sky130_fd_sc_hd__xnor2_2 c404 (.A(net848),
    .B(net823),
    .Y(net358));
 sky130_fd_sc_hd__clkbuf_2 c405 (.A(net831),
    .X(net359));
 sky130_fd_sc_hd__xnor2_2 c406 (.A(net359),
    .B(net356),
    .Y(net360));
 sky130_fd_sc_hd__a21bo_1 c407 (.A1(net360),
    .A2(net356),
    .B1_N(net823),
    .X(net361));
 sky130_fd_sc_hd__xnor2_2 c408 (.A(net353),
    .B(net823),
    .Y(net362));
 sky130_fd_sc_hd__dfrtp_1 c409 (.CLK(clknet_leaf_12_clk),
    .D(net358),
    .RESET_B(net359),
    .Q(net363));
 sky130_fd_sc_hd__dfrtp_1 c410 (.CLK(clknet_leaf_3_clk),
    .D(net356),
    .RESET_B(net358),
    .Q(net364));
 sky130_fd_sc_hd__dfrtp_1 c411 (.CLK(clknet_leaf_3_clk),
    .D(net361),
    .RESET_B(net358),
    .Q(net365));
 sky130_fd_sc_hd__dfsbp_1 c412 (.CLK(clknet_leaf_3_clk),
    .D(net362),
    .SET_B(net360),
    .Q(net366));
 sky130_fd_sc_hd__a21bo_1 c413 (.A1(net351),
    .A2(net357),
    .B1_N(net363),
    .X(net367));
 sky130_fd_sc_hd__a41o_1 c414 (.A1(net357),
    .A2(net360),
    .A3(net359),
    .A4(net823),
    .B1(net338),
    .X(net368));
 sky130_fd_sc_hd__a31o_1 c415 (.A1(net366),
    .A2(net364),
    .A3(net360),
    .B1(net823),
    .X(net369));
 sky130_fd_sc_hd__sdfxbp_1 c416 (.CLK(clknet_leaf_12_clk),
    .D(net863),
    .SCD(net367),
    .SCE(net369),
    .Q(net371),
    .Q_N(net370));
 sky130_fd_sc_hd__sdfxtp_1 c417 (.CLK(clknet_leaf_12_clk),
    .D(net876),
    .SCD(net362),
    .SCE(net358),
    .Q(net372));
 sky130_fd_sc_hd__sdfxtp_1 c418 (.CLK(clknet_leaf_12_clk),
    .D(net861),
    .SCD(net359),
    .SCE(net362),
    .Q(net373));
 sky130_fd_sc_hd__mux4_1 c419 (.A0(net935),
    .A1(net369),
    .A2(net362),
    .A3(net370),
    .S0(net360),
    .S1(net823),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 c420 (.A(net721),
    .X(net375));
 sky130_fd_sc_hd__buf_1 c421 (.A(net264),
    .X(net376));
 sky130_fd_sc_hd__dfsbp_1 c422 (.CLK(clknet_leaf_13_clk),
    .D(net376),
    .SET_B(net823),
    .Q(net378),
    .Q_N(net377));
 sky130_fd_sc_hd__dfstp_2 c423 (.CLK(clknet_leaf_2_clk),
    .D(net376),
    .SET_B(net837),
    .Q(net379));
 sky130_fd_sc_hd__xnor2_4 c424 (.A(net375),
    .B(net379),
    .Y(net380));
 sky130_fd_sc_hd__xnor2_4 c425 (.A(net375),
    .B(net380),
    .Y(net381));
 sky130_fd_sc_hd__xnor2_1 c426 (.A(net379),
    .B(net380),
    .Y(net382));
 sky130_fd_sc_hd__xnor2_1 c427 (.A(net380),
    .B(net931),
    .Y(net383));
 sky130_fd_sc_hd__dfstp_1 c428 (.CLK(clknet_leaf_13_clk),
    .D(net382),
    .SET_B(net383),
    .Q(net384));
 sky130_fd_sc_hd__dfstp_1 c429 (.CLK(clknet_leaf_2_clk),
    .D(net376),
    .SET_B(net381),
    .Q(net385));
 sky130_fd_sc_hd__dlrbn_1 c430 (.D(net898),
    .GATE_N(clknet_leaf_2_clk),
    .RESET_B(net381),
    .Q(net387),
    .Q_N(net386));
 sky130_fd_sc_hd__dlrbn_1 c431 (.D(net387),
    .GATE_N(clknet_leaf_13_clk),
    .RESET_B(net383),
    .Q(net389),
    .Q_N(net388));
 sky130_fd_sc_hd__xnor2_1 c432 (.A(net378),
    .B(net375),
    .Y(net390));
 sky130_fd_sc_hd__sdfxtp_1 c433 (.CLK(clknet_leaf_13_clk),
    .D(net383),
    .SCD(net388),
    .SCE(net380),
    .Q(net391));
 sky130_fd_sc_hd__a21bo_1 c434 (.A1(net917),
    .A2(net389),
    .B1_N(net390),
    .X(net392));
 sky130_fd_sc_hd__dfbbn_1 c435 (.CLK_N(clknet_leaf_13_clk),
    .D(net865),
    .RESET_B(net390),
    .SET_B(net382),
    .Q(net393));
 sky130_fd_sc_hd__dfbbn_1 c436 (.CLK_N(clknet_leaf_13_clk),
    .D(net872),
    .RESET_B(net390),
    .SET_B(net381),
    .Q(net395),
    .Q_N(net394));
 sky130_fd_sc_hd__a21bo_1 c437 (.A1(net380),
    .A2(net393),
    .B1_N(net394),
    .X(net396));
 sky130_fd_sc_hd__dfbbp_1 c438 (.CLK(clknet_leaf_13_clk),
    .D(net392),
    .RESET_B(net396),
    .SET_B(net386),
    .Q(net397));
 sky130_fd_sc_hd__sdfxbp_1 c439 (.CLK(clknet_leaf_13_clk),
    .D(net949),
    .SCD(net395),
    .SCE(net396),
    .Q(net398));
 sky130_fd_sc_hd__sdfxbp_1 c440 (.CLK(clknet_leaf_13_clk),
    .D(net866),
    .SCD(net395),
    .SCE(net392),
    .Q(net399));
 sky130_fd_sc_hd__buf_1 c441 (.A(net696),
    .X(net400));
 sky130_fd_sc_hd__buf_1 c442 (.A(net824),
    .X(net401));
 sky130_fd_sc_hd__xnor2_4 c443 (.A(net938),
    .B(net824),
    .Y(net402));
 sky130_fd_sc_hd__xnor2_1 c444 (.A(net402),
    .B(net401),
    .Y(net403));
 sky130_fd_sc_hd__xnor2_2 c445 (.A(net402),
    .B(net824),
    .Y(net404));
 sky130_fd_sc_hd__a21bo_1 c446 (.A1(net404),
    .A2(net402),
    .B1_N(net824),
    .X(net405));
 sky130_fd_sc_hd__buf_1 c447 (.A(net695),
    .X(net406));
 sky130_fd_sc_hd__xnor2_1 c448 (.A(net824),
    .B(net404),
    .Y(net407));
 sky130_fd_sc_hd__xnor2_1 c449 (.A(net401),
    .B(net406),
    .Y(net408));
 sky130_fd_sc_hd__sdfxtp_1 c450 (.CLK(clknet_leaf_22_clk),
    .D(net402),
    .SCD(net400),
    .SCE(net407),
    .Q(net409));
 sky130_fd_sc_hd__sdfxtp_1 c451 (.CLK(clknet_leaf_28_clk),
    .D(net305),
    .SCD(net405),
    .SCE(net824),
    .Q(net410));
 sky130_fd_sc_hd__xnor2_1 c452 (.A(net409),
    .B(net403),
    .Y(net411));
 sky130_fd_sc_hd__sdfbbn_1 c453 (.CLK_N(clknet_leaf_22_clk),
    .D(net408),
    .RESET_B(net411),
    .SCD(net401),
    .SCE(net402),
    .SET_B(net824),
    .Q(net413),
    .Q_N(net412));
 sky130_fd_sc_hd__xnor2_1 c454 (.A(net946),
    .B(net413),
    .Y(net414));
 sky130_fd_sc_hd__sdfxtp_1 c455 (.CLK(clknet_leaf_22_clk),
    .D(net407),
    .SCD(net414),
    .SCE(net406),
    .Q(net415));
 sky130_fd_sc_hd__a41o_1 c456 (.A1(net413),
    .A2(net415),
    .A3(net409),
    .A4(net824),
    .B1(net408),
    .X(net416));
 sky130_fd_sc_hd__mux4_1 c457 (.A0(net276),
    .A1(net403),
    .A2(net411),
    .A3(net824),
    .S0(net412),
    .S1(net402),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 c458 (.A0(net411),
    .A1(net414),
    .A2(net412),
    .A3(net401),
    .S0(net405),
    .S1(net824),
    .X(net418));
 sky130_fd_sc_hd__sedfxtp_1 c459 (.CLK(clknet_leaf_23_clk),
    .D(net403),
    .DE(net416),
    .SCD(net400),
    .SCE(net926),
    .Q(net419));
 sky130_fd_sc_hd__a21bo_2 c460 (.A1(net404),
    .A2(net840),
    .B1_N(net723),
    .X(net810));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net406),
    .A1(net411),
    .A2(net810),
    .A3(net419),
    .S0(net722),
    .S1(net957),
    .X(net420));
 sky130_fd_sc_hd__buf_1 c462 (.A(net724),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 c463 (.A(net700),
    .X(net421));
 sky130_fd_sc_hd__xnor2_1 c464 (.A(clknet_1_0__leaf_net805),
    .B(net421),
    .Y(net422));
 sky130_fd_sc_hd__xnor2_1 c465 (.A(clknet_1_1__leaf_net805),
    .B(clknet_1_1__leaf_net422),
    .Y(net803));
 sky130_fd_sc_hd__xnor2_1 c466 (.A(net421),
    .B(clknet_1_0__leaf_net805),
    .Y(net423));
 sky130_fd_sc_hd__xnor2_1 c467 (.A(net423),
    .B(clknet_1_0__leaf_net805),
    .Y(net424));
 sky130_fd_sc_hd__clkbuf_2 c468 (.A(net699),
    .X(net425));
 sky130_fd_sc_hd__xnor2_1 c469 (.A(net425),
    .B(clknet_1_0__leaf_net422),
    .Y(net813));
 sky130_fd_sc_hd__xnor2_1 c470 (.A(net425),
    .B(clknet_1_0__leaf_net422),
    .Y(net426));
 sky130_fd_sc_hd__dlrbp_1 c471 (.D(clknet_1_0__leaf_net813),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(clknet_1_1__leaf_net424),
    .Q(net427));
 sky130_fd_sc_hd__mux4_1 c472 (.A0(net427),
    .A1(net425),
    .A2(clknet_1_1__leaf_net805),
    .A3(clknet_1_0__leaf_net803),
    .S0(clknet_1_1__leaf_net422),
    .S1(net421),
    .X(net428));
 sky130_fd_sc_hd__dlrbp_1 c473 (.D(clknet_1_0__leaf_net424),
    .GATE(clknet_leaf_24_clk),
    .RESET_B(clknet_1_0__leaf_net725),
    .Q(net430),
    .Q_N(net429));
 sky130_fd_sc_hd__xnor2_1 c474 (.A(net430),
    .B(net425),
    .Y(net431));
 sky130_fd_sc_hd__xnor2_1 c475 (.A(net421),
    .B(clknet_1_1__leaf_net725),
    .Y(net432));
 sky130_fd_sc_hd__xnor2_1 c476 (.A(clknet_1_0__leaf_net422),
    .B(clknet_1_0__leaf_net725),
    .Y(net433));
 sky130_fd_sc_hd__dlrtn_1 c477 (.D(net431),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(clknet_1_0__leaf_net424),
    .Q(net434));
 sky130_fd_sc_hd__dlrtn_1 c478 (.D(clknet_1_0__leaf_net426),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net432),
    .Q(net435));
 sky130_fd_sc_hd__mux4_1 c479 (.A0(net434),
    .A1(net433),
    .A2(clknet_1_0__leaf_net426),
    .A3(net429),
    .S0(net425),
    .S1(net421),
    .X(net436));
 sky130_fd_sc_hd__dlrtn_1 c480 (.D(clknet_1_0__leaf_net813),
    .GATE_N(clknet_leaf_24_clk),
    .RESET_B(net434),
    .Q(net437));
 sky130_fd_sc_hd__xnor2_1 c481 (.A(net435),
    .B(clknet_1_1__leaf_net726),
    .Y(net808));
 sky130_fd_sc_hd__mux4_1 c482 (.A0(clknet_1_0__leaf_net808),
    .A1(net437),
    .A2(net421),
    .A3(net434),
    .S0(clknet_1_1__leaf_net426),
    .S1(clknet_1_0__leaf_net726),
    .X(net438));
 sky130_fd_sc_hd__buf_4 c504 (.X(net439));
 sky130_fd_sc_hd__xnor2_4 c505 (.A(net439),
    .B(net825),
    .Y(net440));
 sky130_fd_sc_hd__xnor2_4 c506 (.A(net440),
    .B(net915),
    .Y(net441));
 sky130_fd_sc_hd__xnor2_2 c507 (.A(net915),
    .B(net441),
    .Y(net442));
 sky130_fd_sc_hd__clkbuf_1 c508 (.A(net692),
    .X(net443));
 sky130_fd_sc_hd__dlrtp_1 c509 (.D(net352),
    .GATE(clknet_leaf_9_clk),
    .RESET_B(net440),
    .Q(net444));
 sky130_fd_sc_hd__xnor2_4 c510 (.A(net328),
    .B(net441),
    .Y(net445));
 sky130_fd_sc_hd__dfbbn_1 c511 (.CLK_N(clknet_leaf_10_clk),
    .D(net444),
    .RESET_B(net441),
    .SET_B(net445),
    .Q(net447),
    .Q_N(net446));
 sky130_fd_sc_hd__dfbbn_1 c512 (.CLK_N(clknet_leaf_10_clk),
    .D(net444),
    .RESET_B(net884),
    .SET_B(net445),
    .Q(net449),
    .Q_N(net448));
 sky130_fd_sc_hd__xnor2_2 c513 (.A(net447),
    .B(net448),
    .Y(net450));
 sky130_fd_sc_hd__dfbbp_1 c514 (.CLK(clknet_leaf_9_clk),
    .D(net442),
    .RESET_B(net449),
    .SET_B(net445),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__sdfxbp_1 c515 (.CLK(clknet_leaf_10_clk),
    .D(net449),
    .SCD(net445),
    .SCE(net442),
    .Q(net454),
    .Q_N(net453));
 sky130_fd_sc_hd__xnor2_1 c516 (.A(net450),
    .B(net443),
    .Y(net455));
 sky130_fd_sc_hd__a21bo_1 c517 (.A1(net455),
    .A2(net444),
    .B1_N(net451),
    .X(net456));
 sky130_fd_sc_hd__sdfbbn_1 c518 (.CLK_N(clknet_leaf_11_clk),
    .D(net441),
    .RESET_B(net450),
    .SCD(net439),
    .SCE(net456),
    .SET_B(net342),
    .Q(net458),
    .Q_N(net457));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net443),
    .A1(net458),
    .A2(net453),
    .A3(net445),
    .S0(net439),
    .S1(net450),
    .X(net459));
 sky130_fd_sc_hd__sdfxbp_1 c520 (.CLK(clknet_leaf_10_clk),
    .D(net945),
    .SCD(net450),
    .SCE(net727),
    .Q(net461),
    .Q_N(net460));
 sky130_fd_sc_hd__a21bo_1 c521 (.A1(net454),
    .A2(net460),
    .B1_N(net455),
    .X(net462));
 sky130_fd_sc_hd__dlrtp_2 c522 (.D(net462),
    .GATE(clknet_leaf_10_clk),
    .RESET_B(net461),
    .Q(net463));
 sky130_fd_sc_hd__sdfrbp_1 c523 (.CLK(clknet_leaf_10_clk),
    .D(net458),
    .RESET_B(net445),
    .SCD(net462),
    .SCE(net728),
    .Q(net464));
 sky130_fd_sc_hd__sdfbbp_1 c524 (.CLK(clknet_leaf_10_clk),
    .D(net879),
    .RESET_B(net869),
    .SCD(net457),
    .SCE(net940),
    .SET_B(net442),
    .Q(net466),
    .Q_N(net465));
 sky130_fd_sc_hd__xnor2_4 c525 (.A(net466),
    .B(net463),
    .Y(net467));
 sky130_fd_sc_hd__xnor2_4 c526 (.A(net467),
    .B(net721),
    .Y(net468));
 sky130_fd_sc_hd__xnor2_1 c527 (.A(net467),
    .B(net823),
    .Y(net469));
 sky130_fd_sc_hd__dlrtp_1 c528 (.D(net469),
    .GATE(clknet_leaf_11_clk),
    .RESET_B(net463),
    .Q(net470));
 sky130_fd_sc_hd__edfxbp_1 c529 (.CLK(clknet_leaf_11_clk),
    .D(net927),
    .DE(net445),
    .Q(net472),
    .Q_N(net471));
 sky130_fd_sc_hd__edfxtp_1 c530 (.CLK(clknet_leaf_11_clk),
    .D(net469),
    .DE(net947),
    .Q(net473));
 sky130_fd_sc_hd__xnor2_1 c531 (.A(net371),
    .B(net470),
    .Y(net474));
 sky130_fd_sc_hd__xnor2_2 c532 (.A(net354),
    .B(net875),
    .Y(net475));
 sky130_fd_sc_hd__sdlclkp_1 c533 (.CLK(clknet_leaf_12_clk),
    .GATE(net475),
    .SCE(net934),
    .GCLK(net476));
 sky130_fd_sc_hd__xnor2_1 c534 (.A(net472),
    .B(net473),
    .Y(net477));
 sky130_fd_sc_hd__a21bo_1 c535 (.A1(net452),
    .A2(net472),
    .B1_N(net470),
    .X(net478));
 sky130_fd_sc_hd__a21bo_1 c536 (.A1(net478),
    .A2(net474),
    .B1_N(net473),
    .X(net479));
 sky130_fd_sc_hd__sdfxtp_1 c537 (.CLK(clknet_leaf_12_clk),
    .D(net476),
    .SCD(net477),
    .SCE(net475),
    .Q(net480));
 sky130_fd_sc_hd__sdfrbp_1 c538 (.CLK(clknet_leaf_12_clk),
    .D(net368),
    .RESET_B(net475),
    .SCD(net478),
    .SCE(net889),
    .Q(net482),
    .Q_N(net481));
 sky130_fd_sc_hd__a21bo_1 c539 (.A1(net473),
    .A2(net480),
    .B1_N(net481),
    .X(net483));
 sky130_fd_sc_hd__a21bo_1 c540 (.A1(net477),
    .A2(net482),
    .B1_N(net474),
    .X(net484));
 sky130_fd_sc_hd__a21bo_1 c541 (.A1(net484),
    .A2(net948),
    .B1_N(net483),
    .X(net485));
 sky130_fd_sc_hd__sdfxtp_1 c542 (.CLK(clknet_leaf_12_clk),
    .D(net889),
    .SCD(net485),
    .SCE(net927),
    .Q(net486));
 sky130_fd_sc_hd__sdfrtn_1 c543 (.CLK_N(clknet_leaf_11_clk),
    .D(net463),
    .RESET_B(net486),
    .SCD(net475),
    .SCE(net483),
    .Q(net487));
 sky130_fd_sc_hd__a21bo_1 c544 (.A1(net487),
    .A2(net483),
    .B1_N(net486),
    .X(net488));
 sky130_fd_sc_hd__mux4_1 c545 (.A0(net488),
    .A1(net928),
    .A2(net481),
    .A3(net478),
    .S0(net473),
    .S1(net717),
    .X(net489));
 sky130_fd_sc_hd__xnor2_4 c546 (.A(net399),
    .B(net468),
    .Y(net490));
 sky130_fd_sc_hd__buf_1 c547 (.X(net689));
 sky130_fd_sc_hd__buf_1 c548 (.A(net688),
    .X(net492));
 sky130_fd_sc_hd__sdlclkp_2 c549 (.CLK(clknet_leaf_13_clk),
    .GATE(net492),
    .SCE(net490),
    .GCLK(net493));
 sky130_fd_sc_hd__xnor2_1 c550 (.A(net479),
    .B(clknet_1_0__leaf_net493),
    .Y(net494));
 sky130_fd_sc_hd__sdlclkp_4 c551 (.CLK(clknet_leaf_22_clk),
    .GATE(net490),
    .SCE(clknet_1_0__leaf_net494),
    .GCLK(net495));
 sky130_fd_sc_hd__dfrbp_1 c552 (.CLK(clknet_leaf_22_clk),
    .D(clknet_1_0__leaf_net495),
    .RESET_B(clknet_1_0__leaf_net494),
    .Q(net496));
 sky130_fd_sc_hd__dfrbp_1 c553 (.CLK(clknet_leaf_13_clk),
    .D(net490),
    .RESET_B(clknet_1_0__leaf_net493),
    .Q(net498),
    .Q_N(net497));
 sky130_fd_sc_hd__xnor2_1 c554 (.A(net491),
    .B(net498),
    .Y(net499));
 sky130_fd_sc_hd__dfrtn_1 c555 (.CLK_N(clknet_leaf_21_clk),
    .D(net496),
    .RESET_B(net490),
    .Q(net500));
 sky130_fd_sc_hd__dfrtp_4 c556 (.CLK(clknet_leaf_13_clk),
    .D(net871),
    .RESET_B(clknet_1_0__leaf_net494),
    .Q(net501));
 sky130_fd_sc_hd__xnor2_2 c557 (.A(net492),
    .B(net501),
    .Y(net502));
 sky130_fd_sc_hd__a21bo_1 c558 (.A1(net500),
    .A2(net502),
    .B1_N(net498),
    .X(net503));
 sky130_fd_sc_hd__xnor2_1 c559 (.A(net502),
    .B(net501),
    .Y(net504));
 sky130_fd_sc_hd__mux4_1 c560 (.A0(clknet_1_1__leaf_net494),
    .A1(net499),
    .A2(net503),
    .A3(clknet_1_1__leaf_net493),
    .S0(clknet_1_0__leaf_net495),
    .S1(net497),
    .X(net505));
 sky130_fd_sc_hd__xnor2_1 c561 (.A(clknet_1_1__leaf_net495),
    .B(clknet_1_0__leaf_net493),
    .Y(net506));
 sky130_fd_sc_hd__xnor2_1 c562 (.A(net504),
    .B(net503),
    .Y(net507));
 sky130_fd_sc_hd__sdfxtp_1 c563 (.CLK(clknet_leaf_14_clk),
    .D(net506),
    .SCD(net490),
    .SCE(net880),
    .Q(net508));
 sky130_fd_sc_hd__dfbbn_1 c564 (.CLK_N(clknet_leaf_14_clk),
    .D(net507),
    .RESET_B(net508),
    .SET_B(net504),
    .Q(net510),
    .Q_N(net509));
 sky130_fd_sc_hd__a41o_1 c565 (.A1(clknet_1_1__leaf_net493),
    .A2(net509),
    .A3(net497),
    .A4(net502),
    .B1(net729),
    .X(net511));
 sky130_fd_sc_hd__mux4_1 c566 (.A0(net511),
    .A1(net499),
    .A2(net502),
    .A3(net503),
    .S0(clknet_1_1__leaf_net493),
    .S1(clknet_1_1__leaf_net494),
    .X(net512));
 sky130_fd_sc_hd__dfxbp_1 c567 (.CLK(clknet_leaf_21_clk),
    .D(net810),
    .Q(net514),
    .Q_N(net513));
 sky130_fd_sc_hd__dfbbn_2 c568 (.CLK_N(clknet_leaf_21_clk),
    .D(net381),
    .RESET_B(net513),
    .SET_B(net810),
    .Q(net516),
    .Q_N(net515));
 sky130_fd_sc_hd__xnor2_4 c569 (.A(net501),
    .B(net515),
    .Y(net517));
 sky130_fd_sc_hd__xnor2_4 c570 (.A(net517),
    .B(net516),
    .Y(net518));
 sky130_fd_sc_hd__xnor2_2 c571 (.A(net518),
    .B(net516),
    .Y(net519));
 sky130_fd_sc_hd__dfrtp_1 c572 (.CLK(clknet_leaf_21_clk),
    .D(net519),
    .RESET_B(net516),
    .Q(net520));
 sky130_fd_sc_hd__xnor2_4 c573 (.A(net514),
    .B(net518),
    .Y(net802));
 sky130_fd_sc_hd__sdfrtp_1 c574 (.CLK(clknet_leaf_21_clk),
    .D(net802),
    .RESET_B(net830),
    .SCD(net515),
    .SCE(net731),
    .Q(net521));
 sky130_fd_sc_hd__sdfrtp_1 c575 (.CLK(clknet_leaf_21_clk),
    .D(net830),
    .RESET_B(net862),
    .SCD(net932),
    .SCE(net519),
    .Q(net522));
 sky130_fd_sc_hd__xnor2_1 c576 (.A(net516),
    .B(net518),
    .Y(net523));
 sky130_fd_sc_hd__dfrtp_1 c577 (.CLK(clknet_leaf_20_clk),
    .D(net517),
    .RESET_B(net523),
    .Q(net524));
 sky130_fd_sc_hd__dfsbp_1 c578 (.CLK(clknet_leaf_23_clk),
    .D(net523),
    .SET_B(net830),
    .Q(net525));
 sky130_fd_sc_hd__dfsbp_1 c579 (.CLK(clknet_leaf_20_clk),
    .D(net883),
    .SET_B(net519),
    .Q(net527),
    .Q_N(net526));
 sky130_fd_sc_hd__mux4_1 c580 (.A0(net527),
    .A1(net516),
    .A2(net519),
    .A3(net522),
    .S0(net518),
    .S1(net802),
    .X(net528));
 sky130_fd_sc_hd__dfstp_1 c581 (.CLK(clknet_leaf_23_clk),
    .D(net870),
    .SET_B(net523),
    .Q(net529));
 sky130_fd_sc_hd__a21bo_1 c582 (.A1(net902),
    .A2(net960),
    .B1_N(net732),
    .X(net530));
 sky130_fd_sc_hd__dfbbp_1 c583 (.CLK(clknet_leaf_20_clk),
    .D(net530),
    .RESET_B(net951),
    .SET_B(net519),
    .Q(net532),
    .Q_N(net531));
 sky130_fd_sc_hd__xnor2_1 c584 (.A(net532),
    .B(net525),
    .Y(net533));
 sky130_fd_sc_hd__sdfbbn_1 c585 (.CLK_N(clknet_leaf_20_clk),
    .D(net521),
    .RESET_B(net527),
    .SCD(net529),
    .SCE(net531),
    .SET_B(net802),
    .Q(net535),
    .Q_N(net534));
 sky130_fd_sc_hd__sdfbbn_1 c586 (.CLK_N(clknet_leaf_20_clk),
    .D(net533),
    .RESET_B(net529),
    .SCD(net925),
    .SCE(net515),
    .SET_B(net802),
    .Q(net536));
 sky130_fd_sc_hd__mux4_2 c587 (.A0(net535),
    .A1(net536),
    .A2(net521),
    .A3(net515),
    .S0(net522),
    .S1(net518),
    .X(net822));
 sky130_fd_sc_hd__dfstp_1 c588 (.CLK(clknet_leaf_19_clk),
    .D(clknet_1_0__leaf_net803),
    .SET_B(net807),
    .Q(net537));
 sky130_fd_sc_hd__dfstp_2 c589 (.CLK(clknet_leaf_20_clk),
    .D(net894),
    .SET_B(net907),
    .Q(net538));
 sky130_fd_sc_hd__xnor2_1 c590 (.A(net537),
    .B(clknet_1_1__leaf_net808),
    .Y(net539));
 sky130_fd_sc_hd__xnor2_1 c591 (.A(clknet_1_0__leaf_net539),
    .B(net538),
    .Y(net540));
 sky130_fd_sc_hd__xnor2_1 c592 (.A(net538),
    .B(clknet_1_0__leaf_net539),
    .Y(net541));
 sky130_fd_sc_hd__dlrbn_1 c593 (.D(clknet_1_0__leaf_net540),
    .GATE_N(clknet_leaf_18_clk),
    .RESET_B(net894),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__dlrbn_1 c594 (.D(net541),
    .GATE_N(clknet_leaf_19_clk),
    .RESET_B(net912),
    .Q(net811),
    .Q_N(net799));
 sky130_fd_sc_hd__dlrbp_1 c595 (.D(net802),
    .GATE(clknet_leaf_20_clk),
    .RESET_B(clknet_1_1__leaf_net540),
    .Q(net545),
    .Q_N(net544));
 sky130_fd_sc_hd__a21bo_2 c596 (.A1(net545),
    .A2(net542),
    .B1_N(net537),
    .X(net546));
 sky130_fd_sc_hd__xnor2_1 c597 (.A(net538),
    .B(net543),
    .Y(net547));
 sky130_fd_sc_hd__xnor2_2 c598 (.A(net811),
    .B(net546),
    .Y(net548));
 sky130_fd_sc_hd__xnor2_1 c599 (.A(net811),
    .B(net546),
    .Y(net549));
 sky130_fd_sc_hd__xnor2_1 c600 (.A(net548),
    .B(net893),
    .Y(net550));
 sky130_fd_sc_hd__dlrbp_1 c601 (.D(clknet_1_0__leaf_net540),
    .GATE(clknet_leaf_18_clk),
    .RESET_B(net550),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__a41o_1 c602 (.A1(net552),
    .A2(net811),
    .A3(clknet_1_1__leaf_net539),
    .A4(net547),
    .B1(net544),
    .X(net553));
 sky130_fd_sc_hd__xnor2_1 c603 (.A(net547),
    .B(net548),
    .Y(net806));
 sky130_fd_sc_hd__mux4_1 c604 (.A0(clknet_1_0__leaf_net553),
    .A1(net806),
    .A2(net546),
    .A3(clknet_1_1__leaf_net540),
    .S0(net538),
    .S1(net799),
    .X(net554));
 sky130_fd_sc_hd__xnor2_1 c605 (.A(net546),
    .B(net549),
    .Y(net798));
 sky130_fd_sc_hd__mux4_1 c606 (.A0(net543),
    .A1(clknet_1_0__leaf_net553),
    .A2(net548),
    .A3(net799),
    .S0(net552),
    .S1(net801),
    .X(net555));
 sky130_fd_sc_hd__sdfbbp_1 c607 (.CLK(clknet_leaf_19_clk),
    .D(clknet_1_1__leaf_net553),
    .RESET_B(net548),
    .SCD(net911),
    .SCE(clknet_1_1__leaf_net539),
    .SET_B(net834),
    .Q(net556));
 sky130_fd_sc_hd__a21bo_1 c608 (.A1(net537),
    .A2(net556),
    .B1_N(net547),
    .X(net800));
 sky130_fd_sc_hd__mux4_2 c62 (.A0(net788),
    .A1(net773),
    .A2(net780),
    .A3(net782),
    .S0(net785),
    .S1(net790),
    .X(net0));
 sky130_fd_sc_hd__xnor2_1 c63 (.A(net4),
    .B(net784),
    .Y(net1));
 sky130_fd_sc_hd__clkbuf_4 c630 (.A(net452),
    .X(net557));
 sky130_fd_sc_hd__xnor2_4 c631 (.A(net557),
    .B(net465),
    .Y(net558));
 sky130_fd_sc_hd__xnor2_2 c632 (.A(net558),
    .B(net557),
    .Y(net559));
 sky130_fd_sc_hd__clkbuf_2 c633 (.A(net697),
    .X(net560));
 sky130_fd_sc_hd__a21bo_1 c634 (.A1(net560),
    .A2(net557),
    .B1_N(net558),
    .X(net561));
 sky130_fd_sc_hd__a21bo_1 c635 (.A1(net439),
    .A2(net560),
    .B1_N(net558),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 c636 (.A(net697),
    .X(net563));
 sky130_fd_sc_hd__dlrtn_1 c637 (.D(net561),
    .GATE_N(clknet_leaf_10_clk),
    .RESET_B(net558),
    .Q(net564));
 sky130_fd_sc_hd__dlrtn_1 c638 (.D(net559),
    .GATE_N(clknet_leaf_15_clk),
    .RESET_B(net558),
    .Q(net565));
 sky130_fd_sc_hd__xnor2_1 c639 (.A(net338),
    .B(net565),
    .Y(net566));
 sky130_fd_sc_hd__xnor2_2 c64 (.A(net3),
    .B(net783),
    .Y(net2));
 sky130_fd_sc_hd__sdfxbp_1 c640 (.CLK(clknet_leaf_15_clk),
    .D(net558),
    .SCD(net559),
    .SCE(net565),
    .Q(net567));
 sky130_fd_sc_hd__sdfxbp_1 c641 (.CLK(clknet_leaf_10_clk),
    .D(net566),
    .SCD(net560),
    .SCE(net559),
    .Q(net569),
    .Q_N(net568));
 sky130_fd_sc_hd__xnor2_1 c642 (.A(net569),
    .B(net560),
    .Y(net570));
 sky130_fd_sc_hd__sdfbbn_1 c643 (.CLK_N(clknet_leaf_15_clk),
    .D(net560),
    .RESET_B(net570),
    .SCD(net568),
    .SCE(net559),
    .SET_B(net558),
    .Q(net571));
 sky130_fd_sc_hd__xnor2_1 c644 (.A(net567),
    .B(net565),
    .Y(net572));
 sky130_fd_sc_hd__a21bo_1 c645 (.A1(net557),
    .A2(net565),
    .B1_N(net568),
    .X(net573));
 sky130_fd_sc_hd__a41o_1 c646 (.A1(net564),
    .A2(net569),
    .A3(net565),
    .A4(net557),
    .B1(net560),
    .X(net574));
 sky130_fd_sc_hd__a41o_1 c647 (.A1(net572),
    .A2(net574),
    .A3(net560),
    .A4(net568),
    .B1(net557),
    .X(net575));
 sky130_fd_sc_hd__a21bo_1 c648 (.A1(net573),
    .A2(net569),
    .B1_N(net574),
    .X(net576));
 sky130_fd_sc_hd__sdfxtp_1 c649 (.CLK(clknet_leaf_15_clk),
    .D(net576),
    .SCD(net575),
    .SCE(net574),
    .Q(net577));
 sky130_fd_sc_hd__xnor2_4 c65 (.A(net741),
    .B(net791),
    .Y(net3));
 sky130_fd_sc_hd__xnor2_1 c650 (.A(net574),
    .B(net577),
    .Y(net578));
 sky130_fd_sc_hd__buf_1 c651 (.X(net677));
 sky130_fd_sc_hd__buf_1 c652 (.A(net579),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 c653 (.A(net676),
    .X(net581));
 sky130_fd_sc_hd__xnor2_4 c654 (.A(net579),
    .B(net342),
    .Y(net582));
 sky130_fd_sc_hd__xnor2_4 c655 (.A(net582),
    .B(net581),
    .Y(net583));
 sky130_fd_sc_hd__xnor2_4 c656 (.A(net581),
    .B(net582),
    .Y(net584));
 sky130_fd_sc_hd__xnor2_2 c657 (.A(net583),
    .B(net579),
    .Y(net585));
 sky130_fd_sc_hd__xnor2_1 c658 (.A(net563),
    .B(net584),
    .Y(net586));
 sky130_fd_sc_hd__xnor2_2 c659 (.A(net583),
    .B(net580),
    .Y(net587));
 sky130_fd_sc_hd__xnor2_4 c66 (.A(net3),
    .B(net775),
    .Y(net4));
 sky130_fd_sc_hd__dlrtn_1 c660 (.D(net580),
    .GATE_N(clknet_leaf_14_clk),
    .RESET_B(net587),
    .Q(net588));
 sky130_fd_sc_hd__sdfxtp_1 c661 (.CLK(clknet_leaf_14_clk),
    .D(net588),
    .SCD(net587),
    .SCE(net585),
    .Q(net589));
 sky130_fd_sc_hd__sdfrtp_1 c662 (.CLK(clknet_leaf_15_clk),
    .D(net571),
    .RESET_B(net585),
    .SCD(net583),
    .SCE(net579),
    .Q(net590));
 sky130_fd_sc_hd__sdfsbp_1 c663 (.CLK(clknet_leaf_14_clk),
    .D(net445),
    .SCD(net892),
    .SCE(net588),
    .SET_B(net583),
    .Q(net592),
    .Q_N(net591));
 sky130_fd_sc_hd__dlrtp_1 c664 (.D(net587),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net589),
    .Q(net593));
 sky130_fd_sc_hd__sdfxtp_1 c665 (.CLK(clknet_leaf_15_clk),
    .D(net586),
    .SCD(net900),
    .SCE(net583),
    .Q(net594));
 sky130_fd_sc_hd__xnor2_1 c666 (.A(net592),
    .B(net589),
    .Y(net595));
 sky130_fd_sc_hd__dfbbn_1 c667 (.CLK_N(clknet_leaf_14_clk),
    .D(net594),
    .RESET_B(net585),
    .SET_B(net587),
    .Q(net597),
    .Q_N(net596));
 sky130_fd_sc_hd__a21bo_1 c668 (.A1(net468),
    .A2(net593),
    .B1_N(net591),
    .X(net598));
 sky130_fd_sc_hd__a21bo_1 c669 (.A1(net597),
    .A2(net590),
    .B1_N(net594),
    .X(net599));
 sky130_fd_sc_hd__xnor2_1 c67 (.A(net4),
    .B(net2),
    .Y(net5));
 sky130_fd_sc_hd__dfbbn_1 c670 (.CLK_N(clknet_leaf_14_clk),
    .D(net598),
    .RESET_B(net589),
    .SET_B(net930),
    .Q(net600));
 sky130_fd_sc_hd__mux4_1 c671 (.A0(net595),
    .A1(net600),
    .A2(net594),
    .A3(net599),
    .S0(net596),
    .S1(net582),
    .X(net601));
 sky130_fd_sc_hd__buf_2 c672 (.A(net582),
    .X(net602));
 sky130_fd_sc_hd__xnor2_1 c673 (.A(net601),
    .B(net602),
    .Y(net603));
 sky130_fd_sc_hd__buf_2 c674 (.X(net604));
 sky130_fd_sc_hd__xnor2_4 c675 (.A(net584),
    .B(net604),
    .Y(net605));
 sky130_fd_sc_hd__buf_2 c676 (.A(net690),
    .X(net606));
 sky130_fd_sc_hd__xnor2_4 c677 (.A(net602),
    .B(net606),
    .Y(net607));
 sky130_fd_sc_hd__dlrtp_1 c678 (.D(net510),
    .GATE(clknet_leaf_21_clk),
    .RESET_B(net605),
    .Q(net608));
 sky130_fd_sc_hd__dlrtp_1 c679 (.D(net508),
    .GATE(clknet_leaf_14_clk),
    .RESET_B(net607),
    .Q(net609));
 sky130_fd_sc_hd__dfrbp_1 c68 (.CLK(clknet_leaf_34_clk),
    .D(net1),
    .RESET_B(net4),
    .Q(net7),
    .Q_N(net6));
 sky130_fd_sc_hd__edfxbp_1 c680 (.CLK(clknet_leaf_18_clk),
    .D(net846),
    .DE(net605),
    .Q(net611),
    .Q_N(net610));
 sky130_fd_sc_hd__xnor2_1 c681 (.A(net609),
    .B(net604),
    .Y(net612));
 sky130_fd_sc_hd__dfbbp_1 c682 (.CLK(clknet_leaf_14_clk),
    .D(net921),
    .RESET_B(net607),
    .SET_B(net839),
    .Q(net614),
    .Q_N(net613));
 sky130_fd_sc_hd__a21bo_1 c683 (.A1(net614),
    .A2(net604),
    .B1_N(net609),
    .X(net615));
 sky130_fd_sc_hd__xnor2_1 c684 (.A(net604),
    .B(net614),
    .Y(net616));
 sky130_fd_sc_hd__sdfsbp_1 c685 (.CLK(clknet_leaf_14_clk),
    .D(net614),
    .SCD(net605),
    .SCE(net607),
    .SET_B(net846),
    .Q(net617));
 sky130_fd_sc_hd__a21bo_1 c686 (.A1(net608),
    .A2(net610),
    .B1_N(net613),
    .X(net618));
 sky130_fd_sc_hd__xnor2_1 c687 (.A(net616),
    .B(net618),
    .Y(net619));
 sky130_fd_sc_hd__sdfxbp_1 c688 (.CLK(clknet_leaf_21_clk),
    .D(net908),
    .SCD(net612),
    .SCE(net607),
    .Q(net621),
    .Q_N(net620));
 sky130_fd_sc_hd__a21bo_1 c689 (.A1(net612),
    .A2(net618),
    .B1_N(net620),
    .X(net622));
 sky130_fd_sc_hd__dfrbp_1 c69 (.CLK(clknet_leaf_34_clk),
    .D(net794),
    .RESET_B(net1),
    .Q(net9),
    .Q_N(net8));
 sky130_fd_sc_hd__edfxtp_1 c690 (.CLK(clknet_leaf_18_clk),
    .D(net605),
    .DE(net895),
    .Q(net623));
 sky130_fd_sc_hd__sdfbbn_1 c691 (.CLK_N(clknet_leaf_21_clk),
    .D(net622),
    .RESET_B(net623),
    .SCD(net613),
    .SCE(net607),
    .SET_B(net616),
    .Q(net624));
 sky130_fd_sc_hd__mux4_1 c692 (.A0(net624),
    .A1(net619),
    .A2(net604),
    .A3(net609),
    .S0(net605),
    .S1(net606),
    .X(net625));
 sky130_fd_sc_hd__xnor2_2 c693 (.A(net606),
    .B(net734),
    .Y(net626));
 sky130_fd_sc_hd__buf_1 c694 (.A(net685),
    .X(net627));
 sky130_fd_sc_hd__xnor2_1 c695 (.A(net627),
    .B(net734),
    .Y(net628));
 sky130_fd_sc_hd__clkbuf_2 c696 (.A(net684),
    .X(net629));
 sky130_fd_sc_hd__xnor2_2 c697 (.A(net629),
    .B(net734),
    .Y(net630));
 sky130_fd_sc_hd__xnor2_2 c698 (.A(net626),
    .B(net630),
    .Y(net631));
 sky130_fd_sc_hd__sdfxbp_1 c699 (.CLK(clknet_leaf_16_clk),
    .D(net607),
    .SCD(net631),
    .SCE(net629),
    .Q(net633),
    .Q_N(net632));
 sky130_fd_sc_hd__a21bo_1 c70 (.A1(net9),
    .A2(net2),
    .B1_N(net759),
    .X(net10));
 sky130_fd_sc_hd__xnor2_1 c700 (.A(net631),
    .B(net847),
    .Y(net634));
 sky130_fd_sc_hd__a21bo_1 c701 (.A1(net628),
    .A2(net633),
    .B1_N(net630),
    .X(net635));
 sky130_fd_sc_hd__a31o_1 c702 (.A1(net627),
    .A2(net630),
    .A3(net635),
    .B1(net632),
    .X(net636));
 sky130_fd_sc_hd__sdfxtp_1 c703 (.CLK(clknet_leaf_16_clk),
    .D(net603),
    .SCD(net635),
    .SCE(net959),
    .Q(net637));
 sky130_fd_sc_hd__sdfxtp_1 c704 (.CLK(clknet_leaf_16_clk),
    .D(net615),
    .SCD(net885),
    .SCE(net636),
    .Q(net638));
 sky130_fd_sc_hd__a31o_1 c705 (.A1(net638),
    .A2(net635),
    .A3(net629),
    .B1(net632),
    .X(net639));
 sky130_fd_sc_hd__sdfxtp_1 c706 (.CLK(clknet_leaf_16_clk),
    .D(net634),
    .SCD(net888),
    .SCE(net639),
    .Q(net640));
 sky130_fd_sc_hd__dfbbn_1 c707 (.CLK_N(clknet_leaf_16_clk),
    .D(net633),
    .RESET_B(net639),
    .SET_B(net640),
    .Q(net642),
    .Q_N(net641));
 sky130_fd_sc_hd__a21bo_1 c708 (.A1(net630),
    .A2(net637),
    .B1_N(net944),
    .X(net643));
 sky130_fd_sc_hd__sdfbbp_1 c709 (.CLK(clknet_leaf_16_clk),
    .D(net636),
    .RESET_B(net642),
    .SCD(net643),
    .SCE(net639),
    .SET_B(net634),
    .Q(net645),
    .Q_N(net644));
 sky130_fd_sc_hd__mux4_1 c71 (.A0(net10),
    .A1(net8),
    .A2(net2),
    .A3(net4),
    .S0(net778),
    .S1(net6),
    .X(net11));
 sky130_fd_sc_hd__a31o_1 c710 (.A1(net955),
    .A2(net643),
    .A3(net632),
    .B1(net644),
    .X(net646));
 sky130_fd_sc_hd__dfbbn_1 c711 (.CLK_N(clknet_leaf_17_clk),
    .D(net631),
    .RESET_B(net643),
    .SET_B(net646),
    .Q(net648),
    .Q_N(net647));
 sky130_fd_sc_hd__dfbbp_1 c712 (.CLK(clknet_leaf_16_clk),
    .D(net924),
    .RESET_B(net956),
    .SET_B(net847),
    .Q(net649));
 sky130_fd_sc_hd__a21bo_1 c713 (.A1(net611),
    .A2(net649),
    .B1_N(net647),
    .X(net650));
 sky130_fd_sc_hd__xnor2_1 c714 (.A(net800),
    .B(net650),
    .Y(net651));
 sky130_fd_sc_hd__sdlclkp_1 c715 (.CLK(clknet_leaf_18_clk),
    .GATE(net648),
    .SCE(net651),
    .GCLK(net652));
 sky130_fd_sc_hd__sdlclkp_2 c716 (.CLK(clknet_leaf_18_clk),
    .GATE(net651),
    .SCE(clknet_1_0__leaf_net652),
    .GCLK(net653));
 sky130_fd_sc_hd__xnor2_1 c717 (.A(clknet_1_0__leaf_net652),
    .B(clknet_1_0__leaf_net653),
    .Y(net654));
 sky130_fd_sc_hd__xnor2_1 c718 (.A(clknet_1_0__leaf_net653),
    .B(clknet_1_1__leaf_net654),
    .Y(net655));
 sky130_fd_sc_hd__xnor2_1 c719 (.A(clknet_1_0__leaf_net654),
    .B(net650),
    .Y(net656));
 sky130_fd_sc_hd__xnor2_1 c72 (.A(net9),
    .B(net702),
    .Y(net12));
 sky130_fd_sc_hd__xnor2_1 c720 (.A(clknet_1_0__leaf_net654),
    .B(clknet_1_0__leaf_net653),
    .Y(net657));
 sky130_fd_sc_hd__a21bo_1 c721 (.A1(clknet_1_0__leaf_net657),
    .A2(clknet_1_1__leaf_net654),
    .B1_N(clknet_1_0__leaf_net655),
    .X(net658));
 sky130_fd_sc_hd__xnor2_1 c722 (.A(clknet_1_1__leaf_net652),
    .B(clknet_1_0__leaf_net656),
    .Y(net659));
 sky130_fd_sc_hd__sdlclkp_4 c723 (.CLK(clknet_leaf_17_clk),
    .GATE(clknet_1_0__leaf_net655),
    .SCE(clknet_1_0__leaf_net659),
    .GCLK(net660));
 sky130_fd_sc_hd__a21bo_1 c724 (.A1(clknet_1_0__leaf_net657),
    .A2(clknet_1_0__leaf_net655),
    .B1_N(clknet_1_0__leaf_net660),
    .X(net661));
 sky130_fd_sc_hd__sdfxbp_1 c725 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_0__leaf_net658),
    .SCD(clknet_1_1__leaf_net654),
    .SCE(clknet_1_0__leaf_net655),
    .Q(net663),
    .Q_N(net662));
 sky130_fd_sc_hd__sdfxbp_1 c726 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_1__leaf_net660),
    .SCD(net878),
    .SCE(clknet_1_1__leaf_net661),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__sdfbbn_1 c727 (.CLK_N(clknet_leaf_18_clk),
    .D(net651),
    .RESET_B(net662),
    .SCD(clknet_1_0__leaf_net659),
    .SCE(net664),
    .SET_B(clknet_1_1__leaf_net653),
    .Q(net667),
    .Q_N(net666));
 sky130_fd_sc_hd__mux4_1 c728 (.A0(clknet_1_1__leaf_net656),
    .A1(clknet_1_0__leaf_net661),
    .A2(net666),
    .A3(clknet_1_1__leaf_net658),
    .S0(net799),
    .S1(clknet_1_1__leaf_net657),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 c729 (.A0(clknet_1_1__leaf_net653),
    .A1(net667),
    .A2(clknet_1_1__leaf_net657),
    .A3(clknet_1_1__leaf_net655),
    .S0(clknet_1_0__leaf_net660),
    .S1(net735),
    .X(net669));
 sky130_fd_sc_hd__dfbbn_1 c73 (.CLK_N(clknet_leaf_34_clk),
    .D(net4),
    .RESET_B(net1),
    .SET_B(net789),
    .Q(net14),
    .Q_N(net13));
 sky130_fd_sc_hd__mux4_1 c730 (.A0(net665),
    .A1(clknet_1_0__leaf_net658),
    .A2(clknet_1_0__leaf_net669),
    .A3(clknet_1_1__leaf_net657),
    .S0(clknet_1_1__leaf_net653),
    .S1(net736),
    .X(net670));
 sky130_fd_sc_hd__sdfxtp_1 c731 (.CLK(clknet_leaf_17_clk),
    .D(clknet_1_1__leaf_net669),
    .SCD(clknet_1_1__leaf_net659),
    .SCE(net882));
 sky130_fd_sc_hd__xnor2_1 c74 (.A(net12),
    .B(net702),
    .Y(net15));
 sky130_fd_sc_hd__a21bo_1 c75 (.A1(net832),
    .A2(net7),
    .B1_N(net702),
    .X(net16));
 sky130_fd_sc_hd__mux4_1 c76 (.A0(net7),
    .A1(net2),
    .A2(net13),
    .A3(net4),
    .S0(net8),
    .S1(net701),
    .X(net17));
 sky130_fd_sc_hd__a21bo_1 c77 (.A1(net3),
    .A2(net15),
    .B1_N(net701),
    .X(net18));
 sky130_fd_sc_hd__dfrtn_1 c78 (.CLK_N(clknet_leaf_34_clk),
    .D(net5),
    .RESET_B(net16),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 c79 (.CLK(clknet_leaf_33_clk),
    .D(net18),
    .RESET_B(net833),
    .Q(net20));
 sky130_fd_sc_hd__a21bo_1 c80 (.A1(net15),
    .A2(net835),
    .B1_N(net4),
    .X(net21));
 sky130_fd_sc_hd__dfbbn_1 c81 (.CLK_N(clknet_leaf_34_clk),
    .D(net17),
    .RESET_B(net18),
    .SET_B(net787),
    .Q(net22));
 sky130_fd_sc_hd__a21bo_1 c82 (.A1(net2),
    .A2(net22),
    .B1_N(net16),
    .X(net23));
 sky130_fd_sc_hd__sdfrbp_2 c83 (.CLK(clknet_leaf_33_clk),
    .D(net23),
    .RESET_B(net836),
    .SCD(net19),
    .SCE(net835),
    .Q(net25),
    .Q_N(net24));
 sky130_fd_sc_hd__xnor2_4 c84 (.A(net914),
    .B(net19),
    .Y(net26));
 sky130_fd_sc_hd__xnor2_4 c85 (.A(net19),
    .B(net26),
    .Y(net27));
 sky130_fd_sc_hd__xnor2_1 c86 (.A(net26),
    .B(net27),
    .Y(net28));
 sky130_fd_sc_hd__dfrtp_4 c87 (.CLK(clknet_leaf_33_clk),
    .D(net28),
    .RESET_B(net27),
    .Q(net29));
 sky130_fd_sc_hd__xnor2_1 c88 (.A(net27),
    .B(net29),
    .Y(net30));
 sky130_fd_sc_hd__xnor2_1 c89 (.A(net26),
    .B(net849),
    .Y(net31));
 sky130_fd_sc_hd__xnor2_1 c90 (.A(net27),
    .B(net26),
    .Y(net32));
 sky130_fd_sc_hd__dfbbp_1 c91 (.CLK(clknet_leaf_33_clk),
    .D(net28),
    .RESET_B(net31),
    .SET_B(net849),
    .Q(net34),
    .Q_N(net33));
 sky130_fd_sc_hd__dfrtp_1 c92 (.CLK(clknet_leaf_32_clk),
    .D(net32),
    .RESET_B(net850),
    .Q(net35));
 sky130_fd_sc_hd__a21bo_1 c93 (.A1(net31),
    .A2(net778),
    .B1_N(net33),
    .X(net36));
 sky130_fd_sc_hd__xnor2_1 c94 (.A(net34),
    .B(net26),
    .Y(net37));
 sky130_fd_sc_hd__dfsbp_1 c95 (.CLK(clknet_leaf_33_clk),
    .D(net28),
    .SET_B(net37),
    .Q(net38));
 sky130_fd_sc_hd__xnor2_1 c96 (.A(net860),
    .B(net34),
    .Y(net39));
 sky130_fd_sc_hd__dfsbp_1 c97 (.CLK(clknet_leaf_33_clk),
    .D(net39),
    .SET_B(net36),
    .Q(net41),
    .Q_N(net40));
 sky130_fd_sc_hd__sdfxbp_1 c98 (.CLK(clknet_leaf_33_clk),
    .D(net30),
    .SCD(net37),
    .SCE(net936),
    .Q(net42));
 sky130_fd_sc_hd__sdfxbp_1 c99 (.CLK(clknet_leaf_30_clk),
    .D(net920),
    .SCD(net860),
    .SCE(net36),
    .Q(net44),
    .Q_N(net43));
 sky130_fd_sc_hd__sdfstp_1 merge732 (.CLK(clknet_leaf_0_clk),
    .D(net103),
    .SCD(net105),
    .SCE(net765),
    .SET_B(net102),
    .Q(net671));
 sky130_fd_sc_hd__sdfstp_1 merge733 (.CLK(clknet_leaf_3_clk),
    .D(net262),
    .SCD(net263),
    .SCE(net919),
    .SET_B(net265),
    .Q(net672));
 sky130_fd_sc_hd__sdfxtp_1 merge734 (.CLK(clknet_leaf_8_clk),
    .D(net215),
    .SCD(net217),
    .Q(net218));
 sky130_fd_sc_hd__sdfxtp_1 merge735 (.CLK(clknet_leaf_9_clk),
    .D(net355),
    .SCD(net823),
    .SCE(net345),
    .Q(net674));
 sky130_fd_sc_hd__sdfstp_1 merge736 (.CLK(clknet_leaf_6_clk),
    .D(net80),
    .SCD(net87),
    .SCE(net95),
    .SET_B(net874),
    .Q(net675));
 sky130_fd_sc_hd__dfbbn_1 merge737 (.CLK_N(clknet_leaf_11_clk),
    .D(net489),
    .RESET_B(net578),
    .Q(net677),
    .Q_N(net676));
 sky130_fd_sc_hd__sedfxbp_2 merge738 (.CLK(clknet_leaf_26_clk),
    .D(net53),
    .DE(net75),
    .SCD(clknet_1_0__leaf_net199),
    .Q(net195),
    .Q_N(net678));
 sky130_fd_sc_hd__dfbbn_1 merge739 (.CLK_N(clknet_leaf_1_clk),
    .D(net145),
    .RESET_B(net147),
    .Q(net681),
    .Q_N(net680));
 sky130_fd_sc_hd__dfbbp_1 merge740 (.CLK(clknet_leaf_28_clk),
    .D(net169),
    .RESET_B(clknet_1_0__leaf_net307),
    .SET_B(net175),
    .Q(net683),
    .Q_N(net682));
 sky130_fd_sc_hd__sdfxbp_1 merge741 (.CLK(clknet_leaf_16_clk),
    .D(net822),
    .SCD(net626),
    .SCE(net628),
    .Q(net685),
    .Q_N(net684));
 sky130_fd_sc_hd__sedfxbp_1 merge742 (.CLK(clknet_leaf_32_clk),
    .D(net53),
    .DE(net51),
    .SCD(net57),
    .SCE(net916),
    .Q(net687),
    .Q_N(net686));
 sky130_fd_sc_hd__sdfxbp_1 merge743 (.CLK(clknet_leaf_22_clk),
    .D(net490),
    .SCD(net937),
    .Q(net689),
    .Q_N(net688));
 sky130_fd_sc_hd__sedfxtp_4 merge744 (.CLK(clknet_leaf_16_clk),
    .D(net603),
    .DE(net602),
    .SCE(net605),
    .Q(net604));
 sky130_fd_sc_hd__sedfxtp_1 merge745 (.CLK(clknet_leaf_4_clk),
    .DE(net239),
    .SCD(net238),
    .SCE(net237),
    .Q(net240));
 sky130_fd_sc_hd__sedfxtp_4 merge746 (.CLK(clknet_leaf_11_clk),
    .D(net352),
    .DE(net342),
    .SCD(net442),
    .Q(net439));
 sky130_fd_sc_hd__dfrbp_1 merge747 (.CLK(clknet_leaf_8_clk),
    .D(net330),
    .RESET_B(net950),
    .Q(net694),
    .Q_N(net693));
 sky130_fd_sc_hd__sdfrbp_1 merge748 (.CLK(clknet_leaf_22_clk),
    .D(net381),
    .RESET_B(net405),
    .SCD(net404),
    .SCE(net402),
    .Q(net696),
    .Q_N(net695));
 sky130_fd_sc_hd__sdfxtp_1 merge749 (.CLK(clknet_leaf_15_clk),
    .D(net557),
    .SCD(net559),
    .SCE(net562),
    .Q(net697));
 sky130_fd_sc_hd__sdfxtp_1 merge750 (.CLK(clknet_leaf_30_clk),
    .D(net172),
    .SCD(net173),
    .SCE(net175),
    .Q(net698));
 sky130_fd_sc_hd__sdfrbp_1 merge751 (.CLK(clknet_leaf_24_clk),
    .D(clknet_1_0__leaf_net805),
    .RESET_B(net841),
    .SCD(clknet_1_1__leaf_net424),
    .SCE(clknet_1_1__leaf_net422),
    .Q(net700),
    .Q_N(net699));
 sky130_fd_sc_hd__dfxbp_1 s752 (.CLK(clknet_leaf_34_clk),
    .D(net11),
    .Q(net702),
    .Q_N(net701));
 sky130_fd_sc_hd__dfxtp_1 s753 (.CLK(clknet_leaf_5_clk),
    .D(net98),
    .Q(net703));
 sky130_fd_sc_hd__dfxtp_1 s754 (.CLK(clknet_leaf_4_clk),
    .D(net107),
    .Q(net704));
 sky130_fd_sc_hd__dfxtp_1 s755 (.CLK(clknet_leaf_1_clk),
    .D(net122),
    .Q(net705));
 sky130_fd_sc_hd__dlclkp_1 s756 (.CLK(clknet_leaf_29_clk),
    .GATE(net162),
    .GCLK(net706));
 sky130_fd_sc_hd__dlclkp_2 s757 (.CLK(clknet_leaf_29_clk),
    .GATE(net164),
    .GCLK(net707));
 sky130_fd_sc_hd__dlclkp_4 s758 (.CLK(clknet_leaf_26_clk),
    .GATE(net194),
    .GCLK(net708));
 sky130_fd_sc_hd__dlxbn_2 s759 (.D(net202),
    .GATE_N(clknet_leaf_27_clk),
    .Q(net709));
 sky130_fd_sc_hd__dlxbn_1 s760 (.D(net204),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net711),
    .Q_N(net710));
 sky130_fd_sc_hd__dlxbp_1 s761 (.D(net212),
    .GATE(clknet_leaf_25_clk),
    .Q(net713),
    .Q_N(net712));
 sky130_fd_sc_hd__dlxtn_1 s762 (.D(net214),
    .GATE_N(clknet_leaf_25_clk),
    .Q(net812));
 sky130_fd_sc_hd__dlxtn_1 s763 (.D(net232),
    .GATE_N(clknet_leaf_8_clk),
    .Q(net714));
 sky130_fd_sc_hd__dlxtn_1 s764 (.D(net235),
    .GATE_N(clknet_leaf_6_clk),
    .Q(net715));
 sky130_fd_sc_hd__dlxtp_1 s765 (.D(net236),
    .GATE(clknet_leaf_6_clk),
    .Q(net716));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s766 (.D(net255),
    .SLEEP_B(clknet_leaf_3_clk),
    .Q(net717));
 sky130_fd_sc_hd__dfxbp_1 s767 (.CLK(clknet_leaf_6_clk),
    .D(net257),
    .Q(net719),
    .Q_N(net718));
 sky130_fd_sc_hd__dfxbp_1 s768 (.CLK(clknet_leaf_28_clk),
    .D(net327),
    .Q(net720));
 sky130_fd_sc_hd__dfxtp_1 s769 (.CLK(clknet_leaf_12_clk),
    .D(net374),
    .Q(net721));
 sky130_fd_sc_hd__dfxtp_1 s770 (.CLK(clknet_leaf_22_clk),
    .D(net417),
    .Q(net722));
 sky130_fd_sc_hd__dfxtp_1 s771 (.CLK(clknet_leaf_23_clk),
    .D(net418),
    .Q(net723));
 sky130_fd_sc_hd__dlclkp_1 s772 (.CLK(clknet_leaf_23_clk),
    .GATE(net420),
    .GCLK(net724));
 sky130_fd_sc_hd__dlclkp_2 s773 (.CLK(clknet_leaf_24_clk),
    .GATE(net428),
    .GCLK(net725));
 sky130_fd_sc_hd__dlclkp_4 s774 (.CLK(clknet_leaf_24_clk),
    .GATE(net436),
    .GCLK(net726));
 sky130_fd_sc_hd__dlxbn_1 s775 (.D(net438),
    .GATE_N(clknet_leaf_24_clk),
    .Q(net809),
    .Q_N(net807));
 sky130_fd_sc_hd__dlxbn_1 s776 (.D(net459),
    .GATE_N(clknet_leaf_10_clk),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__dlxbp_1 s777 (.D(net505),
    .GATE(clknet_leaf_14_clk),
    .Q(net730),
    .Q_N(net729));
 sky130_fd_sc_hd__dlxtn_1 s778 (.D(net512),
    .GATE_N(clknet_leaf_21_clk),
    .Q(net731));
 sky130_fd_sc_hd__dlxtn_1 s779 (.D(net528),
    .GATE_N(clknet_leaf_20_clk),
    .Q(net732));
 sky130_fd_sc_hd__dlxtn_1 s780 (.D(net554),
    .GATE_N(clknet_leaf_19_clk),
    .Q(net801));
 sky130_fd_sc_hd__dlxtp_1 s781 (.D(net555),
    .GATE(clknet_leaf_19_clk),
    .Q(net733));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s782 (.D(net625),
    .SLEEP_B(clknet_leaf_18_clk),
    .Q(net734));
 sky130_fd_sc_hd__dfxbp_1 s783 (.CLK(clknet_leaf_19_clk),
    .D(net668),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__dfxbp_1 s784 (.CLK(clknet_leaf_17_clk),
    .D(net670),
    .Q(net737));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net679));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in12),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input7 (.A(in14),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in16),
    .X(net745));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net748));
 sky130_fd_sc_hd__buf_1 input13 (.A(in2),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net750));
 sky130_fd_sc_hd__buf_1 input15 (.A(in21),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in22),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(in23),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in24),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input19 (.A(in25),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in26),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in27),
    .X(net757));
 sky130_fd_sc_hd__buf_1 input22 (.A(in28),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in29),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in3),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(in30),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in31),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in33),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in34),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(in35),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in36),
    .X(net766));
 sky130_fd_sc_hd__buf_1 input31 (.A(in37),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in38),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in39),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input34 (.A(in4),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in40),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in41),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in42),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in43),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in44),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(in45),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input41 (.A(in46),
    .X(net777));
 sky130_fd_sc_hd__buf_1 input42 (.A(in47),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(in48),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(in49),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in5),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(in50),
    .X(net782));
 sky130_fd_sc_hd__buf_1 input47 (.A(in51),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net943),
    .X(net784));
 sky130_fd_sc_hd__buf_1 input49 (.A(in53),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(in54),
    .X(net786));
 sky130_fd_sc_hd__buf_1 input51 (.A(in55),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(in56),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(in57),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(in58),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(in59),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(in6),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(in60),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(in61),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in7),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(in8),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(in9),
    .X(net797));
 sky130_fd_sc_hd__buf_2 output62 (.A(net798),
    .X(out10));
 sky130_fd_sc_hd__buf_2 output63 (.A(net799),
    .X(out14));
 sky130_fd_sc_hd__buf_2 output64 (.A(net800),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output65 (.A(net801),
    .X(out17));
 sky130_fd_sc_hd__buf_2 output66 (.A(net802),
    .X(out20));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(clknet_1_1__leaf_net803),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output68 (.A(net804),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(clknet_1_1__leaf_net805),
    .X(out26));
 sky130_fd_sc_hd__buf_2 output70 (.A(net806),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output71 (.A(net807),
    .X(out30));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(clknet_1_0__leaf_net808),
    .X(out33));
 sky130_fd_sc_hd__buf_2 output73 (.A(net809),
    .X(out34));
 sky130_fd_sc_hd__buf_2 output74 (.A(net810),
    .X(out36));
 sky130_fd_sc_hd__buf_2 output75 (.A(net811),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output76 (.A(net812),
    .X(out40));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(clknet_1_1__leaf_net813),
    .X(out41));
 sky130_fd_sc_hd__buf_2 output78 (.A(net814),
    .X(out42));
 sky130_fd_sc_hd__buf_2 output79 (.A(net815),
    .X(out44));
 sky130_fd_sc_hd__buf_2 output80 (.A(net816),
    .X(out45));
 sky130_fd_sc_hd__buf_2 output81 (.A(net817),
    .X(out47));
 sky130_fd_sc_hd__buf_2 output82 (.A(net818),
    .X(out48));
 sky130_fd_sc_hd__buf_6 output83 (.A(clknet_1_0__leaf_net819),
    .X(out50));
 sky130_fd_sc_hd__buf_2 output84 (.A(net820),
    .X(out56));
 sky130_fd_sc_hd__buf_2 output85 (.A(net821),
    .X(out58));
 sky130_fd_sc_hd__buf_2 output86 (.A(net822),
    .X(out7));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(net354),
    .X(net823));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(net400),
    .X(net824));
 sky130_fd_sc_hd__buf_2 max_cap89 (.A(net716),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net195),
    .X(net826));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(net195),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_2 max_cap92 (.A(net245),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net726 (.A(net726),
    .X(clknet_0_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_0__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net726 (.A(clknet_0_net726),
    .X(clknet_1_1__leaf_net726));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net808 (.A(net808),
    .X(clknet_0_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_0__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net808 (.A(clknet_0_net808),
    .X(clknet_1_1__leaf_net808));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net539 (.A(net539),
    .X(clknet_0_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_0__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net539 (.A(clknet_0_net539),
    .X(clknet_1_1__leaf_net539));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net553 (.A(net553),
    .X(clknet_0_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_0__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net553 (.A(clknet_0_net553),
    .X(clknet_1_1__leaf_net553));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net540 (.A(net540),
    .X(clknet_0_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_0__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net540 (.A(clknet_0_net540),
    .X(clknet_1_1__leaf_net540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net725 (.A(net725),
    .X(clknet_0_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_0__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net725 (.A(clknet_0_net725),
    .X(clknet_1_1__leaf_net725));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net805 (.A(net805),
    .X(clknet_0_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_0__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net805 (.A(clknet_0_net805),
    .X(clknet_1_1__leaf_net805));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net424 (.A(net424),
    .X(clknet_0_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_0__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net424 (.A(clknet_0_net424),
    .X(clknet_1_1__leaf_net424));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net803 (.A(net803),
    .X(clknet_0_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_0__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net803 (.A(clknet_0_net803),
    .X(clknet_1_1__leaf_net803));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net422 (.A(net422),
    .X(clknet_0_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_0__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net422 (.A(clknet_0_net422),
    .X(clknet_1_1__leaf_net422));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net426 (.A(net426),
    .X(clknet_0_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_0__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net426 (.A(clknet_0_net426),
    .X(clknet_1_1__leaf_net426));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net813 (.A(net813),
    .X(clknet_0_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_0__leaf_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net813 (.A(clknet_0_net813),
    .X(clknet_1_1__leaf_net813));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net708 (.A(net708),
    .X(clknet_0_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_0__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net708 (.A(clknet_0_net708),
    .X(clknet_1_1__leaf_net708));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net306 (.A(net306),
    .X(clknet_0_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net306 (.A(clknet_0_net306),
    .X(clknet_1_0__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net306 (.A(net829),
    .X(clknet_1_1__leaf_net306));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net316 (.A(net316),
    .X(clknet_0_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_0__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net316 (.A(clknet_0_net316),
    .X(clknet_1_1__leaf_net316));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net819 (.A(net819),
    .X(clknet_0_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_0__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net819 (.A(clknet_0_net819),
    .X(clknet_1_1__leaf_net819));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net198 (.A(net198),
    .X(clknet_0_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_0__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net198 (.A(clknet_0_net198),
    .X(clknet_1_1__leaf_net198));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net200 (.A(net200),
    .X(clknet_0_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_0__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net200 (.A(clknet_0_net200),
    .X(clknet_1_1__leaf_net200));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net199 (.A(net199),
    .X(clknet_0_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_0__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net199 (.A(clknet_0_net199),
    .X(clknet_1_1__leaf_net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net707 (.A(net707),
    .X(clknet_0_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_0__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net707 (.A(clknet_0_net707),
    .X(clknet_1_1__leaf_net707));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net660 (.A(net660),
    .X(clknet_0_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_0__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_1__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net669 (.A(net669),
    .X(clknet_0_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net669 (.A(clknet_0_net669),
    .X(clknet_1_0__leaf_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net669 (.A(clknet_0_net669),
    .X(clknet_1_1__leaf_net669));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net661 (.A(net661),
    .X(clknet_0_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net661 (.A(clknet_0_net661),
    .X(clknet_1_0__leaf_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net661 (.A(clknet_0_net661),
    .X(clknet_1_1__leaf_net661));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net653 (.A(net653),
    .X(clknet_0_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_0__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net653 (.A(clknet_0_net653),
    .X(clknet_1_1__leaf_net653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net658 (.A(net658),
    .X(clknet_0_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_0__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net658 (.A(clknet_0_net658),
    .X(clknet_1_1__leaf_net658));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net654 (.A(net654),
    .X(clknet_0_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_0__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net654 (.A(clknet_0_net654),
    .X(clknet_1_1__leaf_net654));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net656 (.A(net656),
    .X(clknet_0_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_0__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net656 (.A(clknet_0_net656),
    .X(clknet_1_1__leaf_net656));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net659 (.A(net659),
    .X(clknet_0_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_0__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net659 (.A(clknet_0_net659),
    .X(clknet_1_1__leaf_net659));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net652 (.A(net652),
    .X(clknet_0_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_1__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net495 (.A(net495),
    .X(clknet_0_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_0__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net495 (.A(clknet_0_net495),
    .X(clknet_1_1__leaf_net495));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net493 (.A(net493),
    .X(clknet_0_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_0__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net493 (.A(clknet_0_net493),
    .X(clknet_1_1__leaf_net493));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net494 (.A(net494),
    .X(clknet_0_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net494 (.A(clknet_0_net494),
    .X(clknet_1_0__leaf_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net494 (.A(clknet_0_net494),
    .X(clknet_1_1__leaf_net494));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net292 (.A(net292),
    .X(clknet_0_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_0__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net292 (.A(clknet_0_net292),
    .X(clknet_1_1__leaf_net292));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net298 (.A(net298),
    .X(clknet_0_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_0__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net298 (.A(clknet_0_net298),
    .X(clknet_1_1__leaf_net298));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net293 (.A(net293),
    .X(clknet_0_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_0__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net293 (.A(clknet_0_net293),
    .X(clknet_1_1__leaf_net293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net294 (.A(net294),
    .X(clknet_0_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_0__leaf_net294));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net294 (.A(clknet_0_net294),
    .X(clknet_1_1__leaf_net294));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(clknet_0_net306),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net520),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net674),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net14),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net16),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net733),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net20),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net21),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net377),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net671),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net608),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net415),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net810),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net297),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net113),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net120),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net712),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net609),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net633),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net343),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net860),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net31),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net128),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net129),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net705),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net272),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net183),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net184),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net118),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net141),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net142),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net29),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net372),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net517),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net365),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net207),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net387),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net398),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net42),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net253),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net461),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net419),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net384),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net389),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net83),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net89),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net471),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net363),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net687),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net663),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net464),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net730),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net190),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net737),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net522),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net446),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net637),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net322),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net136),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net638),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net480),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net211),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net208),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net590),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net542),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net537),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net621),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net126),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net182),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net385),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net47),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net593),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net220),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net524),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net203),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net137),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net81),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net179),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net802),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net617),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net223),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net72),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net551),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net538),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net189),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net25),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net439),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net58),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net391),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net240),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net251),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net38),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net498),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net268),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net295),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net645),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net534),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net723),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net470),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net487),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net33),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net599),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net379),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net521),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net703),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net473),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net373),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net40),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net282),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net300),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net161),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net463),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net121),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net672),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(in52),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net641),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net456),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net410),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net470),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net482),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net397),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net328),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net529),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net56),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net248),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net693),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net640),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net646),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net723),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net254),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net632),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net526),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net300),
    .X(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in25));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in26));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in27));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in28));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in29));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in30));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(in31));
 sky130_fd_sc_hd__diode_2 ANTENNA_c273_A (.DIODE(in32));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(in33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(in34));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(in35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(in36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(in37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(in38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(in39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(in40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(in41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(in42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(in43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(in44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(in45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(in46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(in47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(in48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(in49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(in50));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(in51));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold115_A (.DIODE(in52));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(in53));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(in54));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(in55));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(in56));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(in57));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(in58));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(in59));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(in60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(in61));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_c639_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c414_B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_S1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c394_B1 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c393_SCD (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c392_A3 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c391_B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_SCE (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_RESET_B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_Q (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge746_DE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c654_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c518_SET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_S0 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_SCE (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_Q_N (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge748_D (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_D (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c436_SET_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c430_RESET_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c429_SET_B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c425_Y (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_c663_D (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c529_DE (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c523_RESET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_A3 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c515_SCD (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c514_SET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c512_SET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_SET_B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_Y (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_s766_Q (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c545_S1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_c294_B (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_X (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_c153_A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold79_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c595_D (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_SET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c585_SET_B (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c580_S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c574_D (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_c573_Y (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_SET_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c567_D (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_A2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_X (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_c356_X (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge741_D (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_c587_X (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
