module netlist_1 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net98;
 wire net99;
 wire net534;
 wire net583;
 wire net731;
 wire net767;
 wire net814;
 wire net864;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net963;
 wire clknet_1_0__leaf_net963;
 wire clknet_1_1__leaf_net963;
 wire clknet_0_net579;
 wire clknet_1_0__leaf_net579;
 wire clknet_1_1__leaf_net579;
 wire clknet_0_net897;
 wire clknet_1_0__leaf_net897;
 wire clknet_1_1__leaf_net897;
 wire clknet_0_net688;
 wire clknet_1_0__leaf_net688;
 wire clknet_1_1__leaf_net688;
 wire clknet_0_net694;
 wire clknet_1_0__leaf_net694;
 wire clknet_1_1__leaf_net694;
 wire clknet_0_net146;
 wire clknet_1_0__leaf_net146;
 wire clknet_1_1__leaf_net146;
 wire clknet_0_net962;
 wire clknet_1_0__leaf_net962;
 wire clknet_1_1__leaf_net962;
 wire clknet_0_net751;
 wire clknet_1_0__leaf_net751;
 wire clknet_1_1__leaf_net751;
 wire clknet_0_net369;
 wire clknet_1_0__leaf_net369;
 wire clknet_1_1__leaf_net369;
 wire clknet_0_net380;
 wire clknet_1_0__leaf_net380;
 wire clknet_1_1__leaf_net380;
 wire clknet_0_net503;
 wire clknet_1_0__leaf_net503;
 wire clknet_1_1__leaf_net503;
 wire clknet_0_net382;
 wire clknet_1_0__leaf_net382;
 wire clknet_1_1__leaf_net382;
 wire clknet_0_net370;
 wire clknet_1_0__leaf_net370;
 wire clknet_1_1__leaf_net370;
 wire clknet_0_net365;
 wire clknet_1_0__leaf_net365;
 wire clknet_1_1__leaf_net365;
 wire clknet_0_net501;
 wire clknet_1_0__leaf_net501;
 wire clknet_1_1__leaf_net501;
 wire clknet_0_net989;
 wire clknet_1_0__leaf_net989;
 wire clknet_1_1__leaf_net989;
 wire clknet_0_net374;
 wire clknet_1_0__leaf_net374;
 wire clknet_1_1__leaf_net374;
 wire clknet_0_net193;
 wire clknet_1_0__leaf_net193;
 wire clknet_1_1__leaf_net193;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net961;
 wire clknet_1_0__leaf_net961;
 wire clknet_1_1__leaf_net961;
 wire clknet_0_net702;
 wire clknet_1_0__leaf_net702;
 wire clknet_1_1__leaf_net702;
 wire clknet_0_net674;
 wire clknet_1_0__leaf_net674;
 wire clknet_1_1__leaf_net674;
 wire clknet_0_net678;
 wire clknet_1_0__leaf_net678;
 wire clknet_1_1__leaf_net678;
 wire clknet_0_net690;
 wire clknet_1_0__leaf_net690;
 wire clknet_1_1__leaf_net690;
 wire clknet_0_net942;
 wire clknet_1_0__leaf_net942;
 wire clknet_1_1__leaf_net942;
 wire clknet_0_net123;
 wire clknet_1_0__leaf_net123;
 wire clknet_1_1__leaf_net123;
 wire clknet_0_net129;
 wire clknet_1_0__leaf_net129;
 wire clknet_1_1__leaf_net129;
 wire clknet_0_net131;
 wire clknet_1_0__leaf_net131;
 wire clknet_1_1__leaf_net131;
 wire clknet_0_net941;
 wire clknet_1_0__leaf_net941;
 wire clknet_1_1__leaf_net941;
 wire clknet_0_net724;
 wire clknet_1_0__leaf_net724;
 wire clknet_1_1__leaf_net724;
 wire clknet_0_net727;
 wire clknet_1_0__leaf_net727;
 wire clknet_1_1__leaf_net727;
 wire clknet_0_net720;
 wire clknet_1_0__leaf_net720;
 wire clknet_1_1__leaf_net720;
 wire clknet_0_net722;
 wire clknet_1_0__leaf_net722;
 wire clknet_1_1__leaf_net722;
 wire clknet_0_net723;
 wire clknet_1_0__leaf_net723;
 wire clknet_1_1__leaf_net723;
 wire clknet_0_net721;
 wire clknet_1_0__leaf_net721;
 wire clknet_1_1__leaf_net721;
 wire clknet_0_net940;
 wire clknet_1_0__leaf_net940;
 wire clknet_1_1__leaf_net940;
 wire clknet_0_net932;
 wire clknet_1_0__leaf_net932;
 wire clknet_1_1__leaf_net932;
 wire clknet_0_net366;
 wire clknet_1_0__leaf_net366;
 wire clknet_1_1__leaf_net366;
 wire clknet_0_net368;
 wire clknet_1_0__leaf_net368;
 wire clknet_1_1__leaf_net368;
 wire clknet_0_net931;
 wire clknet_1_0__leaf_net931;
 wire clknet_1_1__leaf_net931;
 wire clknet_0_net140;
 wire clknet_1_0__leaf_net140;
 wire clknet_1_1__leaf_net140;
 wire clknet_0_net153;
 wire clknet_1_0__leaf_net153;
 wire clknet_1_1__leaf_net153;
 wire clknet_0_net144;
 wire clknet_1_0__leaf_net144;
 wire clknet_1_1__leaf_net144;
 wire clknet_0_net145;
 wire clknet_1_0__leaf_net145;
 wire clknet_1_1__leaf_net145;
 wire clknet_0_net142;
 wire clknet_1_0__leaf_net142;
 wire clknet_1_1__leaf_net142;
 wire clknet_0_net141;
 wire clknet_1_0__leaf_net141;
 wire clknet_1_1__leaf_net141;
 wire clknet_0_net128;
 wire clknet_1_0__leaf_net128;
 wire clknet_1_1__leaf_net128;
 wire clknet_0_net121;
 wire clknet_1_0__leaf_net121;
 wire clknet_1_1__leaf_net121;
 wire clknet_0_net998;
 wire clknet_1_0__leaf_net998;
 wire clknet_1_1__leaf_net998;
 wire clknet_0_net895;
 wire clknet_1_0__leaf_net895;
 wire clknet_1_1__leaf_net895;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;

 sky130_fd_sc_hd__and2_0 c100 (.A(net76),
    .B(net65),
    .X(net77));
 sky130_fd_sc_hd__and2_0 c101 (.A(net74),
    .B(net73),
    .X(net78));
 sky130_fd_sc_hd__and2_1 c102 (.A(net69),
    .B(net65),
    .X(net79));
 sky130_fd_sc_hd__or4bb_1 c103 (.A(net78),
    .B(net79),
    .C_N(net1000),
    .D_N(net71),
    .X(net80));
 sky130_fd_sc_hd__or4bb_1 c104 (.A(net71),
    .B(net1000),
    .C_N(net56),
    .D_N(clknet_1_1__leaf_net895),
    .X(net81));
 sky130_fd_sc_hd__a2111o_1 c105 (.A1(net77),
    .A2(net81),
    .B1(net79),
    .C1(net73),
    .D1(net71),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 c106 (.A(net776),
    .X(net83));
 sky130_fd_sc_hd__and2_0 c107 (.A(net73),
    .B(net83),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 c108 (.A(net790),
    .X(net85));
 sky130_fd_sc_hd__and2_0 c109 (.A(net85),
    .B(net71),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 c110 (.A(net1000),
    .X(net87));
 sky130_fd_sc_hd__buf_1 c111 (.A(net86),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 c112 (.A(net1000),
    .X(net89));
 sky130_fd_sc_hd__and2_2 c113 (.A(net87),
    .B(net89),
    .X(net90));
 sky130_fd_sc_hd__and2_0 c114 (.A(net90),
    .B(net89),
    .X(net91));
 sky130_fd_sc_hd__and2_1 c115 (.A(net90),
    .B(net89),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 c116 (.A(net733),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 c117 (.A(net733),
    .X(net94));
 sky130_fd_sc_hd__and2_0 c118 (.A(net94),
    .B(net89),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 c119 (.A(net831),
    .X(net96));
 sky130_fd_sc_hd__and2_0 c120 (.A(net96),
    .B(net1000),
    .X(net97));
 sky130_fd_sc_hd__and2_1 c121 (.A(net95),
    .B(net90),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 c122 (.A(net1031),
    .X(net99));
 sky130_fd_sc_hd__and2_0 c123 (.A(net93),
    .B(net96),
    .X(net100));
 sky130_fd_sc_hd__and2_0 c124 (.A(net88),
    .B(net97),
    .X(net101));
 sky130_fd_sc_hd__dfbbn_1 c125 (.CLK_N(clknet_4_13_0_clk),
    .D(net99),
    .RESET_B(net92),
    .SET_B(net93),
    .Q(net103),
    .Q_N(net102));
 sky130_fd_sc_hd__clkbuf_1 c126 (.A(net917),
    .X(net104));
 sky130_fd_sc_hd__dfbbp_1 c127 (.CLK(clknet_4_13_0_clk),
    .D(net101),
    .RESET_B(net98),
    .SET_B(net90),
    .Q(net106),
    .Q_N(net105));
 sky130_fd_sc_hd__a2111o_1 c128 (.A1(net97),
    .A2(net104),
    .B1(net105),
    .C1(net102),
    .D1(net95),
    .X(net107));
 sky130_fd_sc_hd__and3_1 c129 (.A(net106),
    .B(net98),
    .C(net107),
    .X(net108));
 sky130_fd_sc_hd__a2111o_1 c130 (.A1(net103),
    .A2(net107),
    .B1(net105),
    .C1(net90),
    .D1(net918),
    .X(net109));
 sky130_fd_sc_hd__sdfxbp_1 c131 (.CLK(clknet_4_13_0_clk),
    .D(net107),
    .SCD(net106),
    .SCE(net1062),
    .Q(net111),
    .Q_N(net110));
 sky130_fd_sc_hd__and2_0 c132 (.A(net814),
    .B(net986),
    .X(net112));
 sky130_fd_sc_hd__and2_2 c133 (.A(net112),
    .B(net985),
    .X(net113));
 sky130_fd_sc_hd__and2_0 c134 (.A(net113),
    .B(net971),
    .X(net114));
 sky130_fd_sc_hd__and2_0 c135 (.A(net112),
    .B(net988),
    .X(net115));
 sky130_fd_sc_hd__and2_2 c136 (.A(net113),
    .B(net974),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 c137 (.A(net879),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 c138 (.A(net879),
    .X(net118));
 sky130_fd_sc_hd__and2_0 c139 (.A(net984),
    .B(net113),
    .X(net119));
 sky130_fd_sc_hd__buf_1 c140 (.A(clknet_1_0__leaf_net931),
    .X(net120));
 sky130_fd_sc_hd__and2_0 c141 (.A(net120),
    .B(net864),
    .X(net121));
 sky130_fd_sc_hd__buf_1 c142 (.A(net773),
    .X(net122));
 sky130_fd_sc_hd__buf_1 c143 (.A(clknet_1_0__leaf_net942),
    .X(net123));
 sky130_fd_sc_hd__and2_1 c144 (.A(net973),
    .B(net122),
    .X(net124));
 sky130_fd_sc_hd__buf_1 c145 (.A(clknet_1_1__leaf_net942),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 c146 (.A(net950),
    .X(net126));
 sky130_fd_sc_hd__or4bb_1 c147 (.A(clknet_1_0__leaf_net123),
    .B(net116),
    .C_N(net126),
    .D_N(net113),
    .X(net127));
 sky130_fd_sc_hd__buf_1 c148 (.A(clknet_1_0__leaf_net931),
    .X(net128));
 sky130_fd_sc_hd__and2_0 c149 (.A(net124),
    .B(clknet_1_1__leaf_net123),
    .X(net129));
 sky130_fd_sc_hd__and2_0 c150 (.A(net113),
    .B(net118),
    .X(net130));
 sky130_fd_sc_hd__and3_1 c151 (.A(clknet_1_0__leaf_net128),
    .B(clknet_1_1__leaf_net129),
    .C(net880),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 c152 (.A0(net117),
    .A1(clknet_1_1__leaf_net131),
    .A2(net130),
    .A3(net116),
    .S0(clknet_1_0__leaf_net128),
    .S1(net113),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 c153 (.A0(net130),
    .A1(clknet_1_0__leaf_net129),
    .A2(clknet_1_1__leaf_net128),
    .A3(clknet_1_0__leaf_net131),
    .S0(net113),
    .S1(net116),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 c154 (.A(net912),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 c155 (.A(net134),
    .X(net135));
 sky130_fd_sc_hd__buf_2 c156 (.A(net135),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 c157 (.A(net764),
    .X(net137));
 sky130_fd_sc_hd__buf_1 c158 (.A(net764),
    .X(net138));
 sky130_fd_sc_hd__and2_2 c159 (.A(net134),
    .B(net936),
    .X(net139));
 sky130_fd_sc_hd__buf_1 c160 (.A(clknet_1_1__leaf_net931),
    .X(net140));
 sky130_fd_sc_hd__and2_0 c161 (.A(net138),
    .B(clknet_1_0__leaf_net140),
    .X(net141));
 sky130_fd_sc_hd__and2_0 c162 (.A(net139),
    .B(clknet_1_0__leaf_net140),
    .X(net142));
 sky130_fd_sc_hd__and3_1 c163 (.A(clknet_1_1__leaf_net141),
    .B(clknet_1_0__leaf_net140),
    .C(net136),
    .X(net143));
 sky130_fd_sc_hd__and2_0 c164 (.A(net134),
    .B(clknet_1_1__leaf_net140),
    .X(net144));
 sky130_fd_sc_hd__and2_0 c165 (.A(clknet_1_0__leaf_net144),
    .B(net878),
    .X(net145));
 sky130_fd_sc_hd__buf_1 c166 (.A(clknet_1_0__leaf_net963),
    .X(net146));
 sky130_fd_sc_hd__and2_0 c167 (.A(clknet_1_0__leaf_net146),
    .B(net138),
    .X(net147));
 sky130_fd_sc_hd__buf_1 c168 (.A(clknet_1_1__leaf_net931),
    .X(net148));
 sky130_fd_sc_hd__and3_1 c169 (.A(net137),
    .B(clknet_1_1__leaf_net142),
    .C(clknet_1_0__leaf_net140),
    .X(net149));
 sky130_fd_sc_hd__and3_1 c170 (.A(net147),
    .B(net148),
    .C(clknet_1_0__leaf_net146),
    .X(net150));
 sky130_fd_sc_hd__sdfxbp_1 c171 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_1__leaf_net145),
    .SCD(clknet_1_1__leaf_net146),
    .SCE(net1054),
    .Q(net152),
    .Q_N(net151));
 sky130_fd_sc_hd__mux4_1 c172 (.A0(clknet_1_0__leaf_net140),
    .A1(clknet_1_0__leaf_net141),
    .A2(net151),
    .A3(net138),
    .S0(net135),
    .S1(net921),
    .X(net153));
 sky130_fd_sc_hd__and3_1 c173 (.A(clknet_1_1__leaf_net153),
    .B(clknet_1_0__leaf_net145),
    .C(clknet_1_1__leaf_net146),
    .X(net154));
 sky130_fd_sc_hd__and3_1 c174 (.A(net150),
    .B(clknet_1_0__leaf_net153),
    .C(net135),
    .X(net155));
 sky130_fd_sc_hd__and3_1 c175 (.A(net136),
    .B(clknet_1_1__leaf_net140),
    .C(net877),
    .X(net156));
 sky130_fd_sc_hd__buf_1 c176 (.A(net35),
    .X(net157));
 sky130_fd_sc_hd__and2_1 c177 (.A(net135),
    .B(net157),
    .X(net158));
 sky130_fd_sc_hd__and2_1 c178 (.A(net35),
    .B(net139),
    .X(net159));
 sky130_fd_sc_hd__buf_1 c179 (.A(net1009),
    .X(net160));
 sky130_fd_sc_hd__and2_0 c180 (.A(net160),
    .B(net152),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 c181 (.A(net747),
    .X(net162));
 sky130_fd_sc_hd__and2_1 c182 (.A(net152),
    .B(net35),
    .X(net163));
 sky130_fd_sc_hd__and2_0 c183 (.A(net161),
    .B(net163),
    .X(net164));
 sky130_fd_sc_hd__and2_1 c184 (.A(net161),
    .B(net163),
    .X(net165));
 sky130_fd_sc_hd__and2_0 c185 (.A(net163),
    .B(net165),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 c186 (.A(net797),
    .X(net167));
 sky130_fd_sc_hd__and2_0 c187 (.A(net162),
    .B(net163),
    .X(net168));
 sky130_fd_sc_hd__or4bb_1 c188 (.A(net159),
    .B(net163),
    .C_N(net168),
    .D_N(net165),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 c189 (.A0(net164),
    .A1(net34),
    .A2(net158),
    .A3(net163),
    .S1(net920),
    .X(net170));
 sky130_fd_sc_hd__and2_0 c190 (.A(net168),
    .B(net888),
    .X(net171));
 sky130_fd_sc_hd__and2_0 c191 (.A(net157),
    .B(net165),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 c192 (.X(net173));
 sky130_fd_sc_hd__clkbuf_1 c193 (.A(net958),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 c194 (.A(net1035),
    .X(net175));
 sky130_fd_sc_hd__a2111o_1 c195 (.A1(net174),
    .A2(net175),
    .B1(net171),
    .C1(net159),
    .D1(net163),
    .X(net176));
 sky130_fd_sc_hd__and2_0 c196 (.A(net165),
    .B(net915),
    .X(net177));
 sky130_fd_sc_hd__sdfxtp_1 c197 (.CLK(clknet_4_7_0_clk),
    .D(net171),
    .SCD(net177),
    .SCE(net914),
    .Q(net178));
 sky130_fd_sc_hd__clkbuf_2 c198 (.A(net178),
    .X(net179));
 sky130_fd_sc_hd__and2_1 c199 (.A(net179),
    .B(net56),
    .X(net180));
 sky130_fd_sc_hd__and2_2 c200 (.A(net62),
    .B(net179),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 c201 (.A(net181),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 c202 (.A(net737),
    .X(net183));
 sky130_fd_sc_hd__buf_1 c203 (.A(net737),
    .X(net184));
 sky130_fd_sc_hd__and2_0 c204 (.A(net179),
    .B(net181),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 c205 (.A(net827),
    .X(net186));
 sky130_fd_sc_hd__buf_1 c206 (.A(net1004),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 c207 (.A(net832),
    .X(net188));
 sky130_fd_sc_hd__and2_1 c208 (.A(net184),
    .B(net186),
    .X(net189));
 sky130_fd_sc_hd__and2_0 c209 (.A(net189),
    .B(net186),
    .X(net190));
 sky130_fd_sc_hd__and3_1 c210 (.A(net187),
    .B(net189),
    .C(net186),
    .X(net191));
 sky130_fd_sc_hd__and3_1 c211 (.A(net188),
    .B(net191),
    .C(net186),
    .X(net192));
 sky130_fd_sc_hd__buf_1 c212 (.A(clknet_1_0__leaf_net962),
    .X(net193));
 sky130_fd_sc_hd__sdfxtp_1 c213 (.CLK(clknet_4_12_0_clk),
    .D(net183),
    .SCD(net192),
    .SCE(net180),
    .Q(net194));
 sky130_fd_sc_hd__mux4_1 c214 (.A0(net194),
    .A1(net190),
    .A2(clknet_1_1__leaf_net193),
    .A3(net189),
    .S0(net191),
    .S1(net179),
    .X(net195));
 sky130_fd_sc_hd__and3_1 c215 (.A(net186),
    .B(clknet_1_0__leaf_net193),
    .C(net191),
    .X(net196));
 sky130_fd_sc_hd__and3_1 c216 (.A(net179),
    .B(net195),
    .C(net194),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 c217 (.A0(clknet_1_1__leaf_net196),
    .A1(net187),
    .A2(net194),
    .A3(net191),
    .S0(net184),
    .X(net198));
 sky130_fd_sc_hd__mux4_1 c218 (.A0(net191),
    .A1(net189),
    .A2(clknet_1_0__leaf_net196),
    .A3(net179),
    .S0(net180),
    .S1(net887),
    .X(net199));
 sky130_fd_sc_hd__sdfxtp_1 c219 (.CLK(clknet_4_13_0_clk),
    .D(net192),
    .SCD(clknet_1_0__leaf_net196),
    .SCE(net1058),
    .Q(net200));
 sky130_fd_sc_hd__and2_1 c220 (.A(net200),
    .B(net56),
    .X(net201));
 sky130_fd_sc_hd__buf_1 c221 (.A(net748),
    .X(net202));
 sky130_fd_sc_hd__buf_1 c222 (.A(net748),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net203),
    .X(net204));
 sky130_fd_sc_hd__and2_1 c224 (.A(net204),
    .B(net1000),
    .X(net205));
 sky130_fd_sc_hd__and2_1 c225 (.A(net84),
    .B(net203),
    .X(net206));
 sky130_fd_sc_hd__and2_1 c226 (.A(net181),
    .B(net205),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 c227 (.A(net791),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 c228 (.A(net823),
    .X(net209));
 sky130_fd_sc_hd__and3_1 c229 (.A(net204),
    .B(net203),
    .C(net208),
    .X(net210));
 sky130_fd_sc_hd__dfbbn_1 c230 (.CLK_N(clknet_4_13_0_clk),
    .D(net206),
    .RESET_B(net210),
    .SET_B(net202),
    .Q(net212),
    .Q_N(net211));
 sky130_fd_sc_hd__or4bb_1 c231 (.A(net212),
    .B(net204),
    .C_N(net210),
    .D_N(net203),
    .X(net213));
 sky130_fd_sc_hd__and3_1 c232 (.A(net205),
    .B(net201),
    .C(net211),
    .X(net214));
 sky130_fd_sc_hd__and3_1 c233 (.A(net209),
    .B(net1000),
    .C(net884),
    .X(net215));
 sky130_fd_sc_hd__and3_1 c234 (.A(net203),
    .B(net210),
    .C(net215),
    .X(net216));
 sky130_fd_sc_hd__and3_1 c235 (.A(net208),
    .B(net207),
    .C(net215),
    .X(net217));
 sky130_fd_sc_hd__and2_1 c236 (.A(net202),
    .B(net205),
    .X(net218));
 sky130_fd_sc_hd__and3_1 c237 (.A(net213),
    .B(net206),
    .C(net212),
    .X(net219));
 sky130_fd_sc_hd__and3_1 c238 (.A(net216),
    .B(net213),
    .C(net916),
    .X(net220));
 sky130_fd_sc_hd__and3_1 c239 (.A(net205),
    .B(net218),
    .C(net883),
    .X(net221));
 sky130_fd_sc_hd__dfbbn_1 c240 (.CLK_N(clknet_4_15_0_clk),
    .D(net218),
    .RESET_B(net911),
    .SET_B(net1015),
    .Q(net223),
    .Q_N(net222));
 sky130_fd_sc_hd__or4bb_1 c241 (.A(net215),
    .B(net223),
    .C_N(net218),
    .D_N(net913),
    .X(net224));
 sky130_fd_sc_hd__and2_0 c242 (.A(net89),
    .B(net915),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 c243 (.A(net225),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 c244 (.A(net759),
    .X(net227));
 sky130_fd_sc_hd__and2_1 c245 (.A(net227),
    .B(net222),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 c246 (.A(net758),
    .X(net229));
 sky130_fd_sc_hd__and2_0 c247 (.A(net89),
    .B(net222),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 c248 (.A(net917),
    .X(net231));
 sky130_fd_sc_hd__and3_1 c249 (.A(net229),
    .B(net1008),
    .C(net231),
    .X(net232));
 sky130_fd_sc_hd__and3_1 c25 (.A(net980),
    .B(net583),
    .C(net976),
    .X(net0));
 sky130_fd_sc_hd__and2_1 c250 (.A(net230),
    .B(net231),
    .X(net233));
 sky130_fd_sc_hd__dfbbp_1 c251 (.CLK(clknet_4_15_0_clk),
    .D(net233),
    .RESET_B(net231),
    .SET_B(net1008),
    .Q(net235),
    .Q_N(net234));
 sky130_fd_sc_hd__and2_0 c252 (.A(net225),
    .B(net231),
    .X(net236));
 sky130_fd_sc_hd__dlymetal6s2s_1 c253 (.A(net842),
    .X(net237));
 sky130_fd_sc_hd__sdfrbp_1 c254 (.CLK(clknet_4_15_0_clk),
    .D(net235),
    .RESET_B(net237),
    .SCD(net233),
    .SCE(net231),
    .Q(net239),
    .Q_N(net238));
 sky130_fd_sc_hd__a2111o_1 c255 (.A1(net237),
    .A2(net236),
    .B1(net228),
    .C1(net231),
    .D1(net1000),
    .X(net240));
 sky130_fd_sc_hd__and3_1 c256 (.A(net235),
    .B(net237),
    .C(net861),
    .X(net241));
 sky130_fd_sc_hd__and2_0 c257 (.A(net241),
    .B(net231),
    .X(net242));
 sky130_fd_sc_hd__and3_1 c258 (.A(net242),
    .B(net1012),
    .C(net237),
    .X(net243));
 sky130_fd_sc_hd__sdfxbp_1 c259 (.CLK(clknet_4_15_0_clk),
    .D(net228),
    .SCD(net242),
    .SCE(net233),
    .Q(net245),
    .Q_N(net244));
 sky130_fd_sc_hd__and2_1 c26 (.A(net0),
    .B(net977),
    .X(net1));
 sky130_fd_sc_hd__and3_1 c260 (.A(net232),
    .B(net1065),
    .C(net1071),
    .X(net246));
 sky130_fd_sc_hd__and3_1 c261 (.A(net243),
    .B(net233),
    .C(net246),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c262 (.A(net246),
    .B(net238),
    .C(net860),
    .X(net248));
 sky130_fd_sc_hd__sdfxbp_1 c263 (.CLK(clknet_4_15_0_clk),
    .D(net248),
    .SCD(net1034),
    .SCE(net237),
    .Q(net250),
    .Q_N(net249));
 sky130_fd_sc_hd__clkbuf_2 c264 (.A(net934),
    .X(net251));
 sky130_fd_sc_hd__and2_1 c265 (.A(net251),
    .B(net936),
    .X(net252));
 sky130_fd_sc_hd__and2_2 c266 (.A(net252),
    .B(net251),
    .X(net253));
 sky130_fd_sc_hd__and2_1 c267 (.A(net251),
    .B(net252),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 c268 (.A(net734),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 c269 (.A(net734),
    .X(net256));
 sky130_fd_sc_hd__and2_1 c27 (.A(net979),
    .B(net1),
    .X(net2));
 sky130_fd_sc_hd__buf_1 c270 (.A(net802),
    .X(net257));
 sky130_fd_sc_hd__and2_1 c271 (.A(net256),
    .B(net251),
    .X(net258));
 sky130_fd_sc_hd__buf_1 c272 (.A(net947),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 c273 (.A(net950),
    .X(net260));
 sky130_fd_sc_hd__and2_0 c274 (.A(net126),
    .B(net258),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 c275 (.A(net773),
    .X(net262));
 sky130_fd_sc_hd__and3_2 c276 (.A(net262),
    .B(net257),
    .C(net258),
    .X(net263));
 sky130_fd_sc_hd__or4bb_1 c277 (.A(net260),
    .B(net263),
    .C_N(net259),
    .D_N(net933),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 c278 (.A(net804),
    .X(net265));
 sky130_fd_sc_hd__buf_1 c279 (.A(net954),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 c28 (.A(net741),
    .X(net3));
 sky130_fd_sc_hd__and3_1 c280 (.A(net255),
    .B(net266),
    .C(net265),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 c281 (.A(net970),
    .X(net268));
 sky130_fd_sc_hd__and3_1 c282 (.A(net259),
    .B(net267),
    .C(net266),
    .X(net269));
 sky130_fd_sc_hd__or4bb_1 c283 (.A(net268),
    .B(net266),
    .C_N(net254),
    .D_N(net265),
    .X(net270));
 sky130_fd_sc_hd__a2111o_1 c284 (.A1(net265),
    .A2(net266),
    .B1(net263),
    .C1(net253),
    .X(net271));
 sky130_fd_sc_hd__mux4_1 c285 (.A0(net269),
    .A1(net259),
    .A2(net265),
    .A3(net253),
    .S0(net863),
    .S1(net934),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 c286 (.A(net922),
    .X(net273));
 sky130_fd_sc_hd__and2_0 c287 (.A(net273),
    .B(net904),
    .X(net274));
 sky130_fd_sc_hd__and2_0 c288 (.A(net273),
    .B(net920),
    .X(net275));
 sky130_fd_sc_hd__and2_1 c289 (.A(net275),
    .B(net273),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c29 (.A(net979),
    .B(net2),
    .C(net987),
    .X(net4));
 sky130_fd_sc_hd__and2_0 c290 (.A(net273),
    .B(net135),
    .X(net277));
 sky130_fd_sc_hd__and3_1 c291 (.A(net273),
    .B(net151),
    .C(net903),
    .X(net278));
 sky130_fd_sc_hd__and2_0 c292 (.A(net278),
    .B(net274),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 c293 (.A(net922),
    .X(net280));
 sky130_fd_sc_hd__and3_1 c294 (.A(net275),
    .B(net280),
    .C(net276),
    .X(net281));
 sky130_fd_sc_hd__and2_0 c295 (.A(net280),
    .B(net278),
    .X(net282));
 sky130_fd_sc_hd__and2_1 c296 (.A(net274),
    .B(net280),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 c297 (.A(net922),
    .X(net284));
 sky130_fd_sc_hd__a2111o_1 c298 (.A1(clknet_1_1__leaf_net144),
    .A2(net283),
    .B1(net281),
    .C1(net253),
    .D1(net273),
    .X(net285));
 sky130_fd_sc_hd__or4bb_1 c299 (.A(net139),
    .B(net284),
    .C_N(net275),
    .D_N(net278),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 c30 (.A(net1011),
    .X(net5));
 sky130_fd_sc_hd__and2_0 c300 (.A(net282),
    .B(net924),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 c301 (.A(net924),
    .X(net288));
 sky130_fd_sc_hd__and3_1 c302 (.A(net283),
    .B(net924),
    .C(net935),
    .X(net289));
 sky130_fd_sc_hd__and3_1 c303 (.A(net289),
    .B(net288),
    .C(net276),
    .X(net290));
 sky130_fd_sc_hd__or4bb_1 c304 (.A(net282),
    .B(net273),
    .C_N(net283),
    .D_N(net1010),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 c305 (.A(net952),
    .X(net292));
 sky130_fd_sc_hd__buf_1 c306 (.A(net812),
    .X(net293));
 sky130_fd_sc_hd__and3_1 c307 (.A(net286),
    .B(net292),
    .C(net291),
    .X(net294));
 sky130_fd_sc_hd__buf_1 c308 (.A(net1018),
    .X(net295));
 sky130_fd_sc_hd__buf_1 c309 (.A(net295),
    .X(net296));
 sky130_fd_sc_hd__and2_0 c31 (.A(net5),
    .B(net767),
    .X(net6));
 sky130_fd_sc_hd__and2_1 c310 (.A(net296),
    .B(net295),
    .X(net297));
 sky130_fd_sc_hd__buf_1 c311 (.A(net1050),
    .X(net298));
 sky130_fd_sc_hd__and2_1 c312 (.A(net298),
    .B(net296),
    .X(net299));
 sky130_fd_sc_hd__and3_2 c313 (.A(net295),
    .B(net298),
    .C(net296),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 c314 (.A(net1050),
    .X(net301));
 sky130_fd_sc_hd__buf_1 c315 (.A(net1067),
    .X(net302));
 sky130_fd_sc_hd__buf_1 c316 (.A(net949),
    .X(net303));
 sky130_fd_sc_hd__and3_1 c317 (.A(net302),
    .B(net303),
    .C(net300),
    .X(net304));
 sky130_fd_sc_hd__and3_1 c318 (.A(net1018),
    .B(net298),
    .C(net303),
    .X(net305));
 sky130_fd_sc_hd__mux4_1 c319 (.A0(net303),
    .A1(net298),
    .A2(net299),
    .A3(net296),
    .S0(net295),
    .S1(net297),
    .X(net306));
 sky130_fd_sc_hd__or4bb_1 c32 (.A(net3),
    .B(net981),
    .C_N(net2),
    .D_N(net1060),
    .X(net7));
 sky130_fd_sc_hd__and3_1 c320 (.A(net303),
    .B(net302),
    .C(net937),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 c321 (.A(net948),
    .X(net308));
 sky130_fd_sc_hd__and3_1 c322 (.A(net305),
    .B(net301),
    .C(net867),
    .X(net309));
 sky130_fd_sc_hd__or4bb_1 c323 (.A(net300),
    .B(net302),
    .C_N(net296),
    .D_N(net1019),
    .X(net310));
 sky130_fd_sc_hd__sdfxtp_1 c324 (.CLK(clknet_4_4_0_clk),
    .D(net158),
    .SCD(net309),
    .SCE(net302),
    .Q(net311));
 sky130_fd_sc_hd__sdfxtp_1 c325 (.CLK(clknet_4_1_0_clk),
    .D(net301),
    .SCD(net297),
    .SCE(net1059),
    .Q(net312));
 sky130_fd_sc_hd__and3_1 c326 (.A(net309),
    .B(net308),
    .C(net312),
    .X(net313));
 sky130_fd_sc_hd__and3_1 c327 (.A(net311),
    .B(net303),
    .C(net937),
    .X(net314));
 sky130_fd_sc_hd__sdfrtn_1 c328 (.CLK_N(clknet_4_4_0_clk),
    .D(net313),
    .RESET_B(net1066),
    .SCD(net296),
    .SCE(net937),
    .Q(net315));
 sky130_fd_sc_hd__mux4_1 c329 (.A0(net308),
    .A1(net293),
    .A2(net297),
    .A3(net311),
    .S0(net867),
    .S1(net937),
    .X(net316));
 sky130_fd_sc_hd__and3_1 c33 (.A(net5),
    .B(net1),
    .C(net2),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 c330 (.A(net762),
    .X(net317));
 sky130_fd_sc_hd__and2_1 c331 (.A(net317),
    .B(net938),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 c332 (.A(net761),
    .X(net319));
 sky130_fd_sc_hd__and2_1 c333 (.A(net319),
    .B(net317),
    .X(net320));
 sky130_fd_sc_hd__and2_1 c334 (.A(net318),
    .B(net181),
    .X(net321));
 sky130_fd_sc_hd__and2_1 c335 (.A(net320),
    .B(net181),
    .X(net322));
 sky130_fd_sc_hd__buf_1 c336 (.A(net817),
    .X(net323));
 sky130_fd_sc_hd__a2111o_1 c337 (.A1(net322),
    .A2(net320),
    .B1(net321),
    .C1(net299),
    .D1(net323),
    .X(net324));
 sky130_fd_sc_hd__and2_0 c338 (.A(net323),
    .B(net317),
    .X(net325));
 sky130_fd_sc_hd__buf_1 c339 (.A(net926),
    .X(net326));
 sky130_fd_sc_hd__and2_2 c34 (.A(net0),
    .B(net6),
    .X(net9));
 sky130_fd_sc_hd__and2_0 c340 (.A(net317),
    .B(net323),
    .X(net327));
 sky130_fd_sc_hd__and2_1 c341 (.A(net327),
    .B(net894),
    .X(net328));
 sky130_fd_sc_hd__and3_1 c342 (.A(net325),
    .B(net326),
    .C(net320),
    .X(net329));
 sky130_fd_sc_hd__a2111o_1 c343 (.A1(net55),
    .A2(net323),
    .B1(net328),
    .C1(net200),
    .D1(net317),
    .X(net330));
 sky130_fd_sc_hd__buf_1 c344 (.A(net819),
    .X(net331));
 sky130_fd_sc_hd__and2_1 c345 (.A(net331),
    .B(net307),
    .X(net332));
 sky130_fd_sc_hd__and2_1 c346 (.A(net312),
    .B(net331),
    .X(net333));
 sky130_fd_sc_hd__mux4_1 c347 (.A0(net299),
    .A1(net329),
    .A2(net333),
    .A3(net320),
    .S0(net332),
    .S1(net317),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 c348 (.A(net952),
    .X(net335));
 sky130_fd_sc_hd__and2_0 c349 (.A(net335),
    .B(net894),
    .X(net336));
 sky130_fd_sc_hd__and3_1 c35 (.A(net3),
    .B(net9),
    .C(net925),
    .X(net10));
 sky130_fd_sc_hd__and2_0 c350 (.A(net326),
    .B(net328),
    .X(net337));
 sky130_fd_sc_hd__mux4_1 c351 (.A0(net337),
    .A1(net335),
    .A2(net333),
    .A3(net322),
    .S0(net320),
    .S1(net181),
    .X(net338));
 sky130_fd_sc_hd__buf_1 c352 (.A(net910),
    .X(net339));
 sky130_fd_sc_hd__buf_1 c353 (.A(net750),
    .X(net340));
 sky130_fd_sc_hd__buf_1 c354 (.A(net340),
    .X(net341));
 sky130_fd_sc_hd__and2_0 c355 (.A(net339),
    .B(net341),
    .X(net342));
 sky130_fd_sc_hd__and2_0 c356 (.A(net342),
    .B(net340),
    .X(net343));
 sky130_fd_sc_hd__and2_0 c357 (.A(net342),
    .B(net341),
    .X(net344));
 sky130_fd_sc_hd__and2_0 c358 (.A(net340),
    .B(net341),
    .X(net345));
 sky130_fd_sc_hd__and3_2 c359 (.A(net341),
    .B(net332),
    .C(net339),
    .X(net346));
 sky130_fd_sc_hd__dfbbn_1 c36 (.CLK_N(clknet_4_4_0_clk),
    .D(net978),
    .RESET_B(net10),
    .SET_B(net9),
    .Q(net12),
    .Q_N(net11));
 sky130_fd_sc_hd__clkbuf_1 c360 (.A(net910),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 c361 (.A(net750),
    .X(net348));
 sky130_fd_sc_hd__and2_1 c362 (.A(net339),
    .B(net341),
    .X(net349));
 sky130_fd_sc_hd__and2_1 c363 (.A(net347),
    .B(net349),
    .X(net350));
 sky130_fd_sc_hd__or4bb_1 c364 (.A(net307),
    .B(net350),
    .C_N(net349),
    .D_N(net1000),
    .X(net351));
 sky130_fd_sc_hd__sdfbbn_1 c365 (.CLK_N(clknet_4_12_0_clk),
    .D(net350),
    .RESET_B(net349),
    .SCD(net341),
    .SCE(net340),
    .SET_B(clknet_1_0__leaf_net932),
    .Q(net353),
    .Q_N(net352));
 sky130_fd_sc_hd__and3_1 c366 (.A(net350),
    .B(net348),
    .C(net342),
    .X(net354));
 sky130_fd_sc_hd__or4bb_1 c367 (.A(net353),
    .B(net344),
    .C_N(net349),
    .D_N(net350),
    .X(net355));
 sky130_fd_sc_hd__or4bb_1 c368 (.A(net345),
    .B(net347),
    .C_N(net352),
    .D_N(net341),
    .X(net356));
 sky130_fd_sc_hd__and2_0 c369 (.A(net349),
    .B(clknet_1_0__leaf_net932),
    .X(net357));
 sky130_fd_sc_hd__or4bb_1 c37 (.A(net9),
    .B(net12),
    .C_N(net731),
    .D_N(net0),
    .X(net13));
 sky130_fd_sc_hd__sdfxtp_1 c370 (.CLK(clknet_4_12_0_clk),
    .D(net356),
    .SCD(net353),
    .SCE(net350),
    .Q(net358));
 sky130_fd_sc_hd__clkbuf_1 c371 (.A(net803),
    .X(net359));
 sky130_fd_sc_hd__dfbbn_1 c372 (.CLK_N(clknet_4_12_0_clk),
    .D(net358),
    .RESET_B(net359),
    .SET_B(net350),
    .Q(net361),
    .Q_N(net360));
 sky130_fd_sc_hd__mux4_1 c373 (.A0(net348),
    .A1(net360),
    .A2(net358),
    .A3(net350),
    .S0(net349),
    .S1(net352),
    .X(net362));
 sky130_fd_sc_hd__and2_1 c374 (.A(net239),
    .B(net110),
    .X(net363));
 sky130_fd_sc_hd__and2_0 c375 (.A(net363),
    .B(net250),
    .X(net364));
 sky130_fd_sc_hd__buf_1 c376 (.A(clknet_1_0__leaf_net751),
    .X(net365));
 sky130_fd_sc_hd__buf_1 c377 (.A(clknet_1_1__leaf_net932),
    .X(net366));
 sky130_fd_sc_hd__and2_1 c378 (.A(net250),
    .B(net363),
    .X(net367));
 sky130_fd_sc_hd__and2_0 c379 (.A(net367),
    .B(clknet_1_0__leaf_net366),
    .X(net368));
 sky130_fd_sc_hd__or4bb_1 c38 (.A(net980),
    .B(net13),
    .C_N(net982),
    .D_N(net9),
    .X(net14));
 sky130_fd_sc_hd__buf_1 c380 (.A(clknet_1_1__leaf_net751),
    .X(net369));
 sky130_fd_sc_hd__and2_0 c381 (.A(net364),
    .B(clknet_1_1__leaf_net369),
    .X(net370));
 sky130_fd_sc_hd__buf_1 c382 (.A(net806),
    .X(net371));
 sky130_fd_sc_hd__and3_1 c383 (.A(clknet_1_0__leaf_net369),
    .B(clknet_1_1__leaf_net368),
    .C(net371),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 c384 (.A(net827),
    .X(net373));
 sky130_fd_sc_hd__and2_0 c385 (.A(clknet_1_1__leaf_net365),
    .B(net866),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 c386 (.A(net826),
    .X(net375));
 sky130_fd_sc_hd__buf_1 c387 (.A(net819),
    .X(net376));
 sky130_fd_sc_hd__dfbbn_1 c388 (.CLK_N(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net374),
    .RESET_B(net367),
    .SET_B(net346),
    .Q(net378),
    .Q_N(net377));
 sky130_fd_sc_hd__and2_0 c389 (.A(net378),
    .B(clknet_1_1__leaf_net369),
    .X(net379));
 sky130_fd_sc_hd__or4bb_1 c39 (.A(net972),
    .B(net9),
    .C_N(net6),
    .D_N(net1024),
    .X(net15));
 sky130_fd_sc_hd__a2111o_1 c390 (.A1(net363),
    .A2(clknet_1_1__leaf_net365),
    .B1(clknet_1_0__leaf_net369),
    .C1(net377),
    .D1(net376),
    .X(net380));
 sky130_fd_sc_hd__and3_1 c391 (.A(net375),
    .B(clknet_1_0__leaf_net374),
    .C(clknet_1_0__leaf_net380),
    .X(net381));
 sky130_fd_sc_hd__a2111o_1 c392 (.A1(clknet_1_1__leaf_net366),
    .A2(net378),
    .B1(clknet_1_1__leaf_net374),
    .C1(clknet_1_1__leaf_net380),
    .D1(clknet_1_1__leaf_net365),
    .X(net382));
 sky130_fd_sc_hd__or4bb_1 c393 (.A(clknet_1_0__leaf_net382),
    .B(net377),
    .C_N(net371),
    .D_N(clknet_1_0__leaf_net374),
    .X(net383));
 sky130_fd_sc_hd__a2111o_1 c394 (.A1(net376),
    .A2(net379),
    .B1(clknet_1_1__leaf_net366),
    .C1(clknet_1_0__leaf_net382),
    .D1(clknet_1_1__leaf_net374),
    .X(net384));
 sky130_fd_sc_hd__a2111o_1 c395 (.A1(clknet_1_1__leaf_net380),
    .A2(net367),
    .B1(clknet_1_1__leaf_net382),
    .C1(net866),
    .D1(net913),
    .X(net385));
 sky130_fd_sc_hd__buf_1 c396 (.A(net928),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 c397 (.A(net386),
    .X(net387));
 sky130_fd_sc_hd__buf_1 c398 (.A(net736),
    .X(net388));
 sky130_fd_sc_hd__and2_1 c399 (.A(net387),
    .B(net388),
    .X(net389));
 sky130_fd_sc_hd__or4bb_1 c40 (.A(net1),
    .B(net15),
    .C_N(net11),
    .D_N(net9),
    .X(net16));
 sky130_fd_sc_hd__and2_0 c400 (.A(net386),
    .B(net388),
    .X(net390));
 sky130_fd_sc_hd__dfbbp_1 c401 (.CLK(clknet_4_0_0_clk),
    .D(net389),
    .RESET_B(net387),
    .SET_B(net253),
    .Q(net392),
    .Q_N(net391));
 sky130_fd_sc_hd__and2_1 c402 (.A(net1027),
    .B(net390),
    .X(net393));
 sky130_fd_sc_hd__sdfrtp_1 c403 (.CLK(clknet_4_0_0_clk),
    .D(net392),
    .RESET_B(net393),
    .SCD(net388),
    .SCE(net387),
    .Q(net394));
 sky130_fd_sc_hd__and2_1 c404 (.A(net394),
    .B(net387),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 c405 (.A(net964),
    .X(net396));
 sky130_fd_sc_hd__sdfxbp_1 c406 (.CLK(clknet_4_0_0_clk),
    .D(net387),
    .SCD(net1051),
    .SCE(net395),
    .Q(net398),
    .Q_N(net397));
 sky130_fd_sc_hd__clkbuf_1 c407 (.A(net735),
    .X(net399));
 sky130_fd_sc_hd__and2_1 c408 (.A(net398),
    .B(net396),
    .X(net400));
 sky130_fd_sc_hd__and2_1 c409 (.A(net122),
    .B(net397),
    .X(net401));
 sky130_fd_sc_hd__or4bb_1 c41 (.A(net6),
    .B(net10),
    .C_N(net3),
    .D_N(net9),
    .X(net17));
 sky130_fd_sc_hd__sdfxbp_1 c410 (.CLK(clknet_4_2_0_clk),
    .D(net389),
    .SCD(net1046),
    .SCE(net400),
    .Q(net403),
    .Q_N(net402));
 sky130_fd_sc_hd__and3_1 c411 (.A(net401),
    .B(net395),
    .C(net402),
    .X(net404));
 sky130_fd_sc_hd__and3_1 c412 (.A(net1068),
    .B(net401),
    .C(net889),
    .X(net405));
 sky130_fd_sc_hd__and3_1 c413 (.A(net405),
    .B(net396),
    .C(net400),
    .X(net406));
 sky130_fd_sc_hd__and3_1 c414 (.A(net393),
    .B(net399),
    .C(net406),
    .X(net407));
 sky130_fd_sc_hd__and3_1 c415 (.A(net406),
    .B(net401),
    .C(net889),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 c416 (.A0(net400),
    .A1(net405),
    .A2(net406),
    .A3(net401),
    .S0(net389),
    .S1(net903),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 c417 (.A0(net388),
    .A1(net1046),
    .A2(net400),
    .A3(net405),
    .S0(net387),
    .S1(net1017),
    .X(net410));
 sky130_fd_sc_hd__buf_1 c418 (.A(net757),
    .X(net411));
 sky130_fd_sc_hd__buf_1 c419 (.A(net411),
    .X(net412));
 sky130_fd_sc_hd__and3_1 c42 (.A(net12),
    .B(net9),
    .C(net925),
    .X(net18));
 sky130_fd_sc_hd__and2_1 c420 (.A(net293),
    .B(net411),
    .X(net413));
 sky130_fd_sc_hd__and2_1 c421 (.A(net413),
    .B(net412),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net412),
    .X(net415));
 sky130_fd_sc_hd__buf_1 c423 (.A(net414),
    .X(net416));
 sky130_fd_sc_hd__and3_1 c424 (.A(net411),
    .B(net413),
    .C(net892),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 c425 (.A(net757),
    .X(net418));
 sky130_fd_sc_hd__and2_1 c426 (.A(net412),
    .B(net415),
    .X(net419));
 sky130_fd_sc_hd__buf_1 c427 (.A(net1069),
    .X(net420));
 sky130_fd_sc_hd__and2_0 c428 (.A(net411),
    .B(net420),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 c429 (.A(net811),
    .X(net422));
 sky130_fd_sc_hd__mux4_2 c43 (.A0(net13),
    .A1(net18),
    .A2(net9),
    .A3(net2),
    .S0(net904),
    .S1(net925),
    .X(net19));
 sky130_fd_sc_hd__and2_0 c430 (.A(net420),
    .B(net421),
    .X(net423));
 sky130_fd_sc_hd__and2_0 c431 (.A(net414),
    .B(net421),
    .X(net424));
 sky130_fd_sc_hd__and3_1 c432 (.A(net417),
    .B(net423),
    .C(net421),
    .X(net425));
 sky130_fd_sc_hd__sdfxtp_1 c433 (.CLK(clknet_4_2_0_clk),
    .D(net418),
    .SCD(net424),
    .SCE(net412),
    .Q(net426));
 sky130_fd_sc_hd__and3_1 c434 (.A(net1005),
    .B(net414),
    .C(net420),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 c435 (.A(net970),
    .X(net428));
 sky130_fd_sc_hd__and3_1 c436 (.A(net423),
    .B(net424),
    .C(net414),
    .X(net429));
 sky130_fd_sc_hd__and2_0 c437 (.A(net1005),
    .B(net1016),
    .X(net430));
 sky130_fd_sc_hd__a2111o_1 c438 (.A1(net430),
    .A2(net422),
    .B1(net428),
    .C1(net1005),
    .D1(net414),
    .X(net431));
 sky130_fd_sc_hd__and3_1 c439 (.A(net287),
    .B(net427),
    .C(net430),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 c44 (.A(net42),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 c440 (.A(net732),
    .X(net433));
 sky130_fd_sc_hd__buf_1 c441 (.A(net314),
    .X(net434));
 sky130_fd_sc_hd__and2_0 c442 (.A(net434),
    .B(net312),
    .X(net435));
 sky130_fd_sc_hd__and2_1 c443 (.A(net434),
    .B(net34),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 c444 (.A(net732),
    .X(net437));
 sky130_fd_sc_hd__and2_2 c445 (.A(net437),
    .B(net434),
    .X(net438));
 sky130_fd_sc_hd__buf_1 c446 (.A(net779),
    .X(net439));
 sky130_fd_sc_hd__and2_0 c447 (.A(net428),
    .B(net437),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 c448 (.A(net793),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 c449 (.A(net1056),
    .X(net442));
 sky130_fd_sc_hd__buf_1 c45 (.A(net42),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 c450 (.A(net800),
    .X(net443));
 sky130_fd_sc_hd__and2_0 c451 (.A(net443),
    .B(net442),
    .X(net444));
 sky130_fd_sc_hd__and2_0 c452 (.A(net315),
    .B(net444),
    .X(net445));
 sky130_fd_sc_hd__and2_2 c453 (.A(net444),
    .B(net442),
    .X(net446));
 sky130_fd_sc_hd__and3_1 c454 (.A(net445),
    .B(net439),
    .C(net442),
    .X(net447));
 sky130_fd_sc_hd__and3_1 c455 (.A(net442),
    .B(net446),
    .C(net438),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 c456 (.A(net812),
    .X(net449));
 sky130_fd_sc_hd__and2_0 c457 (.A(net440),
    .B(net434),
    .X(net450));
 sky130_fd_sc_hd__sdfbbn_1 c458 (.CLK_N(clknet_4_9_0_clk),
    .D(net449),
    .RESET_B(net446),
    .SCD(net438),
    .SCE(net442),
    .SET_B(net876),
    .Q(net452),
    .Q_N(net451));
 sky130_fd_sc_hd__buf_6 c459 (.A(net944),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 c46 (.A(net21),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 c460 (.A0(net436),
    .A1(net450),
    .A2(net452),
    .A3(net453),
    .S0(net446),
    .S1(net442),
    .X(net454));
 sky130_fd_sc_hd__sdfbbp_1 c461 (.CLK(clknet_4_9_0_clk),
    .D(net442),
    .RESET_B(net453),
    .SCD(net446),
    .SCE(net438),
    .SET_B(net1032),
    .Q(net456),
    .Q_N(net455));
 sky130_fd_sc_hd__and2_0 c462 (.A(net456),
    .B(net332),
    .X(net457));
 sky130_fd_sc_hd__and2_2 c463 (.A(net336),
    .B(net318),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 c464 (.A(net332),
    .X(net459));
 sky130_fd_sc_hd__buf_2 c465 (.A(net458),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 c466 (.A(net760),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_2 c467 (.A(net760),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 c468 (.A(net794),
    .X(net463));
 sky130_fd_sc_hd__and2_2 c469 (.A(net319),
    .B(net462),
    .X(net464));
 sky130_fd_sc_hd__and2_1 c47 (.A(net986),
    .B(net1024),
    .X(net23));
 sky130_fd_sc_hd__and3_1 c470 (.A(net463),
    .B(net462),
    .C(net464),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 c471 (.A(net794),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 c472 (.A(net946),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 c473 (.A(net818),
    .X(net468));
 sky130_fd_sc_hd__and2_0 c474 (.A(net461),
    .B(net464),
    .X(net469));
 sky130_fd_sc_hd__and3_2 c475 (.A(net465),
    .B(net466),
    .C(net455),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 c476 (.A(net960),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 c477 (.A(net849),
    .X(net472));
 sky130_fd_sc_hd__mux4_1 c478 (.A0(net467),
    .A1(net471),
    .A2(net464),
    .A3(net470),
    .S0(net460),
    .S1(net462),
    .X(net473));
 sky130_fd_sc_hd__sdfxtp_1 c479 (.CLK(clknet_4_12_0_clk),
    .D(net318),
    .SCD(net462),
    .SCE(net470),
    .Q(net474));
 sky130_fd_sc_hd__clkbuf_1 c48 (.A(net743),
    .X(net24));
 sky130_fd_sc_hd__buf_1 c480 (.A(net811),
    .X(net475));
 sky130_fd_sc_hd__mux4_1 c481 (.A0(net474),
    .A1(net469),
    .A2(net475),
    .A3(net458),
    .S0(net462),
    .S1(net461),
    .X(net476));
 sky130_fd_sc_hd__buf_2 c482 (.A(net779),
    .X(net477));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net475),
    .A1(net477),
    .A2(net470),
    .A3(net474),
    .S0(net464),
    .S1(net460),
    .X(net478));
 sky130_fd_sc_hd__and3_1 c484 (.A(net477),
    .B(net181),
    .C(net923),
    .X(net479));
 sky130_fd_sc_hd__dlymetal6s2s_1 c485 (.A(net765),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 c486 (.A(net765),
    .X(net481));
 sky130_fd_sc_hd__and2_1 c487 (.A(net361),
    .B(net480),
    .X(net482));
 sky130_fd_sc_hd__and2_0 c488 (.A(net482),
    .B(net480),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 c489 (.A(net483),
    .X(net994));
 sky130_fd_sc_hd__buf_1 c49 (.A(net23),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 c490 (.A(net1045),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 c491 (.A(net1052),
    .X(net485));
 sky130_fd_sc_hd__and3_1 c492 (.A(net481),
    .B(net482),
    .C(net484),
    .X(net486));
 sky130_fd_sc_hd__and2_1 c493 (.A(net480),
    .B(net483),
    .X(net487));
 sky130_fd_sc_hd__buf_1 c494 (.A(net821),
    .X(net488));
 sky130_fd_sc_hd__and3_2 c495 (.A(net483),
    .B(net484),
    .C(net477),
    .X(net489));
 sky130_fd_sc_hd__and3_1 c496 (.A(net485),
    .B(net486),
    .C(net480),
    .X(net490));
 sky130_fd_sc_hd__buf_1 c497 (.A(net945),
    .X(net491));
 sky130_fd_sc_hd__buf_1 c498 (.A(net816),
    .X(net492));
 sky130_fd_sc_hd__and3_1 c499 (.A(net486),
    .B(net492),
    .C(net480),
    .X(net493));
 sky130_fd_sc_hd__and2_0 c50 (.A(net20),
    .B(net21),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c500 (.A(net484),
    .B(net492),
    .X(net494));
 sky130_fd_sc_hd__mux4_1 c501 (.A0(net490),
    .A1(net486),
    .A2(net484),
    .A3(net489),
    .S0(net477),
    .S1(net491),
    .X(net495));
 sky130_fd_sc_hd__and3_1 c502 (.A(net494),
    .B(net490),
    .C(net926),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 c503 (.A(net926),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 c504 (.A(net810),
    .X(net498));
 sky130_fd_sc_hd__a2111o_1 c505 (.A1(net488),
    .A2(net492),
    .B1(net498),
    .C1(net480),
    .D1(net484),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 c509 (.A(net744),
    .X(net500));
 sky130_fd_sc_hd__and2_2 c51 (.A(net24),
    .B(net25),
    .X(net27));
 sky130_fd_sc_hd__and2_0 c510 (.A(clknet_1_1__leaf_net365),
    .B(net923),
    .X(net501));
 sky130_fd_sc_hd__and2_0 c511 (.A(clknet_1_0__leaf_net365),
    .B(net911),
    .X(net502));
 sky130_fd_sc_hd__and2_0 c512 (.A(clknet_1_0__leaf_net380),
    .B(net249),
    .X(net503));
 sky130_fd_sc_hd__dlymetal6s2s_1 c513 (.A(net744),
    .X(net996));
 sky130_fd_sc_hd__buf_1 c514 (.A(net795),
    .X(net504));
 sky130_fd_sc_hd__buf_1 c515 (.A(net966),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 c516 (.A(net803),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_1 c517 (.A(net960),
    .X(net506));
 sky130_fd_sc_hd__or4bb_1 c518 (.A(net506),
    .B(net505),
    .C_N(clknet_1_1__leaf_net501),
    .D_N(net996),
    .X(net989));
 sky130_fd_sc_hd__mux4_1 c519 (.A0(net497),
    .A1(clknet_1_0__leaf_net989),
    .A2(net996),
    .A3(net504),
    .S0(clknet_1_0__leaf_net503),
    .S1(clknet_1_0__leaf_net365),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_1 c52 (.A(net743),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 c520 (.A(net951),
    .X(net508));
 sky130_fd_sc_hd__or4bb_1 c521 (.A(net502),
    .B(net505),
    .C_N(clknet_1_1__leaf_net503),
    .D_N(clknet_1_0__leaf_net501),
    .X(net509));
 sky130_fd_sc_hd__and2_0 c522 (.A(net373),
    .B(net504),
    .X(net510));
 sky130_fd_sc_hd__and2_4 c523 (.A(net504),
    .B(net505),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 c524 (.A(net956),
    .X(net991));
 sky130_fd_sc_hd__mux4_1 c525 (.A0(net508),
    .A1(net250),
    .A2(net511),
    .A3(net505),
    .S0(clknet_1_1__leaf_net365),
    .S1(net902),
    .X(net512));
 sky130_fd_sc_hd__and2_1 c526 (.A(net510),
    .B(net511),
    .X(net993));
 sky130_fd_sc_hd__or4bb_4 c527 (.A(clknet_1_1__leaf_net365),
    .B(net512),
    .C_N(net511),
    .D_N(net902),
    .X(net999));
 sky130_fd_sc_hd__buf_1 c528 (.A(net745),
    .X(net513));
 sky130_fd_sc_hd__buf_1 c529 (.A(net513),
    .X(net514));
 sky130_fd_sc_hd__buf_1 c53 (.A(net854),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 c530 (.A(net745),
    .X(net515));
 sky130_fd_sc_hd__and2_0 c531 (.A(net514),
    .B(net513),
    .X(net516));
 sky130_fd_sc_hd__and2_0 c532 (.A(net515),
    .B(net513),
    .X(net517));
 sky130_fd_sc_hd__and2_0 c533 (.A(net517),
    .B(net513),
    .X(net518));
 sky130_fd_sc_hd__buf_1 c534 (.A(net518),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 c535 (.A(net799),
    .X(net520));
 sky130_fd_sc_hd__and2_1 c536 (.A(net518),
    .B(net520),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_1 c537 (.A(net796),
    .X(net522));
 sky130_fd_sc_hd__sdfxtp_1 c538 (.CLK(clknet_4_2_0_clk),
    .D(net516),
    .SCD(net519),
    .SCE(net515),
    .Q(net523));
 sky130_fd_sc_hd__clkbuf_1 c539 (.A(net798),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_2 c54 (.A(net1026),
    .X(net30));
 sky130_fd_sc_hd__and2_0 c540 (.A(net524),
    .B(net522),
    .X(net525));
 sky130_fd_sc_hd__and2_1 c541 (.A(net525),
    .B(net522),
    .X(net526));
 sky130_fd_sc_hd__and2_0 c542 (.A(net517),
    .B(net525),
    .X(net527));
 sky130_fd_sc_hd__and2_0 c543 (.A(net520),
    .B(net526),
    .X(net528));
 sky130_fd_sc_hd__and2_0 c544 (.A(net527),
    .B(net526),
    .X(net529));
 sky130_fd_sc_hd__or4bb_1 c545 (.A(net526),
    .B(net527),
    .C_N(net523),
    .D_N(net529),
    .X(net530));
 sky130_fd_sc_hd__dfbbn_1 c546 (.CLK_N(clknet_4_8_0_clk),
    .D(net528),
    .RESET_B(net529),
    .SET_B(net526),
    .Q(net532),
    .Q_N(net531));
 sky130_fd_sc_hd__and3_1 c547 (.A(net529),
    .B(net532),
    .C(net526),
    .X(net533));
 sky130_fd_sc_hd__and2_0 c548 (.A(net528),
    .X(net927));
 sky130_fd_sc_hd__dfbbn_1 c549 (.CLK_N(clknet_4_8_0_clk),
    .D(net521),
    .RESET_B(net526),
    .SET_B(net927),
    .Q(net536),
    .Q_N(net535));
 sky130_fd_sc_hd__clkbuf_1 c55 (.A(net953),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 c550 (.A(net536),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 c551 (.A(net537),
    .X(net538));
 sky130_fd_sc_hd__buf_1 c552 (.A(net537),
    .X(net539));
 sky130_fd_sc_hd__and2_0 c553 (.A(net537),
    .B(net539),
    .X(net540));
 sky130_fd_sc_hd__and2_2 c554 (.A(net539),
    .B(net538),
    .X(net541));
 sky130_fd_sc_hd__dfbbp_1 c555 (.CLK(clknet_4_2_0_clk),
    .D(net540),
    .RESET_B(net538),
    .SET_B(net537),
    .Q(net543),
    .Q_N(net542));
 sky130_fd_sc_hd__and2_1 c556 (.A(net415),
    .B(net537),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 c557 (.A(net738),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 c558 (.A(net1028),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 c559 (.A(net796),
    .X(net547));
 sky130_fd_sc_hd__and2_1 c56 (.A(net21),
    .B(net30),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 c560 (.A(net807),
    .X(net548));
 sky130_fd_sc_hd__and3_1 c561 (.A(net541),
    .B(net537),
    .C(net539),
    .X(net549));
 sky130_fd_sc_hd__and2_0 c562 (.A(net545),
    .B(net537),
    .X(net550));
 sky130_fd_sc_hd__buf_1 c563 (.A(net802),
    .X(net551));
 sky130_fd_sc_hd__and3_1 c564 (.A(net547),
    .B(net550),
    .C(net551),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 c565 (.A(net959),
    .X(net553));
 sky130_fd_sc_hd__and2_0 c566 (.A(net551),
    .B(net547),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c567 (.A(net552),
    .B(net554),
    .C(net551),
    .X(net555));
 sky130_fd_sc_hd__and3_1 c568 (.A(net538),
    .B(net551),
    .C(net885),
    .X(net556));
 sky130_fd_sc_hd__and3_1 c569 (.A(net539),
    .B(net553),
    .C(net531),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_1 c57 (.A(net1064),
    .X(net33));
 sky130_fd_sc_hd__sdfbbn_1 c570 (.CLK_N(clknet_4_8_0_clk),
    .D(net548),
    .RESET_B(net552),
    .SCD(net557),
    .SCE(net537),
    .SET_B(net539),
    .Q(net559),
    .Q_N(net558));
 sky130_fd_sc_hd__and3_1 c571 (.A(net546),
    .B(net558),
    .C(net556),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 c572 (.A(net869),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 c573 (.A(net938),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 c574 (.A(net905),
    .X(net563));
 sky130_fd_sc_hd__and2_1 c575 (.A(net550),
    .B(net453),
    .X(net564));
 sky130_fd_sc_hd__and3_4 c576 (.A(net453),
    .B(net562),
    .C(net561),
    .X(net565));
 sky130_fd_sc_hd__and2_0 c577 (.A(net561),
    .B(net456),
    .X(net566));
 sky130_fd_sc_hd__and2_0 c578 (.A(net563),
    .B(net561),
    .X(net567));
 sky130_fd_sc_hd__and2_4 c579 (.A(net565),
    .B(net561),
    .X(net568));
 sky130_fd_sc_hd__sdfrbp_2 c58 (.CLK(clknet_4_5_0_clk),
    .D(net33),
    .RESET_B(net32),
    .SCD(net28),
    .SCE(net30),
    .Q(net35),
    .Q_N(net34));
 sky130_fd_sc_hd__clkbuf_1 c580 (.A(net742),
    .X(net569));
 sky130_fd_sc_hd__and2_0 c581 (.A(net567),
    .B(net561),
    .X(net570));
 sky130_fd_sc_hd__and2_0 c582 (.A(net453),
    .B(net561),
    .X(net571));
 sky130_fd_sc_hd__sdfxbp_1 c583 (.CLK(clknet_4_9_0_clk),
    .D(net566),
    .SCD(net568),
    .SCE(net564),
    .Q(net573),
    .Q_N(net572));
 sky130_fd_sc_hd__clkbuf_1 c584 (.A(net742),
    .X(net574));
 sky130_fd_sc_hd__and2_0 c585 (.A(net569),
    .B(net571),
    .X(net575));
 sky130_fd_sc_hd__and2_1 c586 (.A(net562),
    .B(net574),
    .X(net576));
 sky130_fd_sc_hd__and2_0 c587 (.A(net576),
    .B(net561),
    .X(net577));
 sky130_fd_sc_hd__buf_1 c588 (.A(net774),
    .X(net578));
 sky130_fd_sc_hd__buf_1 c589 (.A(clknet_1_1__leaf_net963),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 c59 (.A(net1047),
    .X(net36));
 sky130_fd_sc_hd__and3_1 c590 (.A(net573),
    .B(clknet_1_1__leaf_net579),
    .C(net576),
    .X(net580));
 sky130_fd_sc_hd__a2111o_1 c591 (.A1(clknet_1_0__leaf_net579),
    .A2(net580),
    .B1(net565),
    .C1(net576),
    .D1(net561),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 c592 (.A(net922),
    .X(net582));
 sky130_fd_sc_hd__mux4_2 c593 (.A0(net582),
    .A1(net576),
    .A2(net573),
    .A3(net568),
    .S0(net565),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_1 c594 (.A(net746),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 c595 (.A(net1022),
    .X(net585));
 sky130_fd_sc_hd__and2_0 c596 (.A(net584),
    .B(net585),
    .X(net586));
 sky130_fd_sc_hd__and2_1 c597 (.A(net585),
    .B(net586),
    .X(net587));
 sky130_fd_sc_hd__sdfxbp_1 c598 (.CLK(clknet_4_9_0_clk),
    .D(net586),
    .SCD(net587),
    .SCE(net477),
    .Q(net589),
    .Q_N(net588));
 sky130_fd_sc_hd__and2_1 c599 (.A(net1022),
    .B(net477),
    .X(net590));
 sky130_fd_sc_hd__and3_1 c60 (.A(net28),
    .B(net35),
    .C(net30),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 c600 (.A(net955),
    .X(net591));
 sky130_fd_sc_hd__and3_1 c601 (.A(net590),
    .B(net589),
    .C(net591),
    .X(net592));
 sky130_fd_sc_hd__and3_2 c602 (.A(net472),
    .B(net592),
    .C(net1070),
    .X(net593));
 sky130_fd_sc_hd__and3_1 c603 (.A(net587),
    .B(net591),
    .C(net585),
    .X(net594));
 sky130_fd_sc_hd__or4bb_1 c604 (.A(net593),
    .B(net585),
    .C_N(net590),
    .D_N(net1002),
    .X(net595));
 sky130_fd_sc_hd__buf_1 c605 (.A(net746),
    .X(net596));
 sky130_fd_sc_hd__sdfxtp_2 c606 (.CLK(clknet_4_11_0_clk),
    .D(net593),
    .SCD(clknet_1_0__leaf_net998),
    .SCE(net899),
    .Q(net597));
 sky130_fd_sc_hd__mux4_1 c607 (.A0(net596),
    .A1(net592),
    .A2(net589),
    .A3(net593),
    .S0(net587),
    .S1(net597),
    .X(net598));
 sky130_fd_sc_hd__sdfxtp_1 c608 (.CLK(clknet_4_11_0_clk),
    .D(net1039),
    .SCD(net1057),
    .SCE(net593),
    .Q(net599));
 sky130_fd_sc_hd__and3_1 c609 (.A(net592),
    .B(net585),
    .C(net1013),
    .X(net600));
 sky130_fd_sc_hd__or4bb_1 c61 (.A(net37),
    .B(net23),
    .C_N(net27),
    .D_N(net30),
    .X(net38));
 sky130_fd_sc_hd__sdfrtp_1 c610 (.CLK(clknet_4_11_0_clk),
    .D(net1042),
    .RESET_B(net1002),
    .SCD(net587),
    .SCE(net939),
    .Q(net601));
 sky130_fd_sc_hd__and3_1 c611 (.A(net599),
    .B(net596),
    .C(net900),
    .X(net602));
 sky130_fd_sc_hd__or4bb_1 c612 (.A(net601),
    .B(net597),
    .C_N(net596),
    .D_N(net591),
    .X(net603));
 sky130_fd_sc_hd__or4bb_1 c613 (.A(net477),
    .B(net597),
    .C_N(net900),
    .D_N(net939),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 c614 (.A0(net602),
    .A1(net604),
    .A2(net601),
    .A3(net599),
    .S0(net585),
    .S1(net588),
    .X(net605));
 sky130_fd_sc_hd__mux4_2 c615 (.A0(net603),
    .A1(net605),
    .A2(net597),
    .A3(net588),
    .S0(net899),
    .S1(net939),
    .X(net606));
 sky130_fd_sc_hd__buf_1 c616 (.A(net769),
    .X(net607));
 sky130_fd_sc_hd__and2_1 c617 (.A(net223),
    .B(net607),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 c618 (.A(net768),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 c619 (.A(net787),
    .X(net610));
 sky130_fd_sc_hd__or4bb_1 c62 (.A(net36),
    .B(net29),
    .C_N(net35),
    .D_N(net871),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 c620 (.A(net607),
    .X(net611));
 sky130_fd_sc_hd__and2_0 c621 (.A(net609),
    .B(net610),
    .X(net612));
 sky130_fd_sc_hd__buf_1 c622 (.A(net609),
    .X(net613));
 sky130_fd_sc_hd__and2_0 c623 (.A(net613),
    .B(net612),
    .X(net614));
 sky130_fd_sc_hd__and3_1 c624 (.A(net611),
    .B(net608),
    .C(net612),
    .X(net615));
 sky130_fd_sc_hd__and2_0 c625 (.A(net612),
    .B(net613),
    .X(net616));
 sky130_fd_sc_hd__and2_2 c626 (.A(net597),
    .B(net615),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_1 c627 (.A(net1038),
    .X(net617));
 sky130_fd_sc_hd__and3_1 c628 (.A(net614),
    .B(net610),
    .C(net997),
    .X(net618));
 sky130_fd_sc_hd__and2_0 c629 (.A(net616),
    .B(net908),
    .X(net619));
 sky130_fd_sc_hd__or4bb_1 c63 (.A(net1048),
    .B(net29),
    .C_N(net27),
    .D_N(net28),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 c630 (.A(net770),
    .X(net620));
 sky130_fd_sc_hd__and2_0 c631 (.A(net610),
    .B(net615),
    .X(net621));
 sky130_fd_sc_hd__a2111o_1 c632 (.A1(net620),
    .A2(net614),
    .B1(net606),
    .C1(net997),
    .D1(net607),
    .X(net622));
 sky130_fd_sc_hd__and3_1 c633 (.A(net346),
    .B(net617),
    .C(net619),
    .X(net623));
 sky130_fd_sc_hd__sdfxtp_1 c634 (.CLK(clknet_4_11_0_clk),
    .D(net615),
    .SCD(net621),
    .SCE(net1043),
    .Q(net992));
 sky130_fd_sc_hd__a2111o_1 c635 (.A1(net621),
    .A2(net608),
    .B1(net620),
    .C1(net997),
    .X(net624));
 sky130_fd_sc_hd__and2_0 c636 (.A(net617),
    .B(net907),
    .X(net625));
 sky130_fd_sc_hd__sdfbbn_1 c637 (.CLK_N(clknet_4_11_0_clk),
    .D(net625),
    .RESET_B(net997),
    .SCD(net607),
    .SCE(net873),
    .SET_B(net907),
    .Q(net990),
    .Q_N(net626));
 sky130_fd_sc_hd__and3_1 c64 (.A(net1053),
    .B(net30),
    .C(net1020),
    .X(net41));
 sky130_fd_sc_hd__buf_1 c65 (.A(in20),
    .X(net42));
 sky130_fd_sc_hd__and2_1 c66 (.A(net41),
    .B(net34),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 c660 (.A(net536),
    .X(net627));
 sky130_fd_sc_hd__buf_1 c661 (.A(net627),
    .X(net628));
 sky130_fd_sc_hd__and2_1 c662 (.A(net628),
    .B(net627),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_1 c663 (.X(net630));
 sky130_fd_sc_hd__and2_0 c664 (.A(net532),
    .B(net627),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 c665 (.A(net766),
    .X(net632));
 sky130_fd_sc_hd__and3_1 c666 (.A(net631),
    .B(net628),
    .C(net627),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 c667 (.A(net820),
    .X(net634));
 sky130_fd_sc_hd__buf_1 c668 (.A(net825),
    .X(net635));
 sky130_fd_sc_hd__and2_1 c669 (.A(net630),
    .B(net628),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 c67 (.A(net43),
    .X(net44));
 sky130_fd_sc_hd__and2_0 c670 (.A(net627),
    .B(net628),
    .X(net637));
 sky130_fd_sc_hd__dfbbn_1 c671 (.CLK_N(clknet_4_8_0_clk),
    .D(net636),
    .RESET_B(net637),
    .SET_B(net633),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__dfbbn_1 c672 (.CLK_N(clknet_4_8_0_clk),
    .D(net637),
    .RESET_B(net636),
    .SET_B(net635),
    .Q(net641),
    .Q_N(net640));
 sky130_fd_sc_hd__sdfbbp_1 c673 (.CLK(clknet_4_10_0_clk),
    .D(net641),
    .RESET_B(net628),
    .SCD(net635),
    .SCE(net636),
    .SET_B(net629),
    .Q(net643),
    .Q_N(net642));
 sky130_fd_sc_hd__and2_0 c674 (.A(net634),
    .B(net639),
    .X(net644));
 sky130_fd_sc_hd__and3_1 c675 (.A(net1063),
    .B(net638),
    .C(net637),
    .X(net645));
 sky130_fd_sc_hd__dfbbp_1 c676 (.CLK(clknet_4_8_0_clk),
    .D(net644),
    .RESET_B(net1063),
    .SET_B(net636),
    .Q(net647),
    .Q_N(net646));
 sky130_fd_sc_hd__and3_1 c677 (.A(net639),
    .B(net642),
    .C(net647),
    .X(net648));
 sky130_fd_sc_hd__a2111o_1 c678 (.A1(net640),
    .A2(net627),
    .B1(net646),
    .C1(net635),
    .D1(net874),
    .X(net649));
 sky130_fd_sc_hd__and3_1 c679 (.A(net648),
    .B(net649),
    .C(net647),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 c68 (.A(net753),
    .X(net45));
 sky130_fd_sc_hd__a2111o_1 c680 (.A1(net635),
    .A2(net649),
    .B1(net638),
    .C1(net627),
    .D1(net631),
    .X(net651));
 sky130_fd_sc_hd__and3_1 c681 (.A(net650),
    .B(net651),
    .C(net1025),
    .X(net652));
 sky130_fd_sc_hd__buf_1 c682 (.A(net647),
    .X(net653));
 sky130_fd_sc_hd__and2_1 c683 (.A(net653),
    .B(net646),
    .X(net654));
 sky130_fd_sc_hd__and2_0 c684 (.A(net654),
    .B(net653),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 c685 (.X(net656));
 sky130_fd_sc_hd__and2_1 c686 (.A(net653),
    .B(net1030),
    .X(net657));
 sky130_fd_sc_hd__and2_1 c687 (.A(net657),
    .B(net654),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_1 c688 (.A(net730),
    .X(net659));
 sky130_fd_sc_hd__and2_0 c689 (.A(net656),
    .B(net654),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 c69 (.A(net45),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 c690 (.A(net808),
    .X(net661));
 sky130_fd_sc_hd__and2_1 c691 (.A(net657),
    .B(net659),
    .X(net662));
 sky130_fd_sc_hd__buf_1 c692 (.A(net820),
    .X(net663));
 sky130_fd_sc_hd__buf_1 c693 (.A(net822),
    .X(net664));
 sky130_fd_sc_hd__and3_1 c694 (.A(net559),
    .B(net654),
    .C(net663),
    .X(net665));
 sky130_fd_sc_hd__and3_1 c695 (.A(net655),
    .B(net659),
    .C(net664),
    .X(net666));
 sky130_fd_sc_hd__and2_1 c696 (.A(net661),
    .B(net891),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_1 c697 (.A(net809),
    .X(net668));
 sky130_fd_sc_hd__mux4_1 c698 (.A0(net659),
    .A1(net663),
    .A2(net664),
    .A3(net657),
    .S0(net665),
    .S1(net653),
    .X(net669));
 sky130_fd_sc_hd__and3_1 c699 (.A(net668),
    .B(net667),
    .C(net653),
    .X(net670));
 sky130_fd_sc_hd__buf_1 c70 (.A(net1021),
    .X(net47));
 sky130_fd_sc_hd__and3_1 c700 (.A(net654),
    .B(net663),
    .C(net891),
    .X(net671));
 sky130_fd_sc_hd__mux4_1 c701 (.A0(net663),
    .A1(net670),
    .A2(net665),
    .A3(net664),
    .S0(net671),
    .S1(net654),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_1 c702 (.A(net943),
    .X(net673));
 sky130_fd_sc_hd__buf_1 c703 (.A(clknet_1_0__leaf_net961),
    .X(net674));
 sky130_fd_sc_hd__buf_1 c704 (.A(net749),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net667),
    .X(net676));
 sky130_fd_sc_hd__buf_1 c706 (.A(net891),
    .X(net677));
 sky130_fd_sc_hd__and2_0 c707 (.A(clknet_1_0__leaf_net674),
    .B(net677),
    .X(net678));
 sky130_fd_sc_hd__and2_0 c708 (.A(net676),
    .B(net677),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 c709 (.A(net749),
    .X(net680));
 sky130_fd_sc_hd__buf_1 c71 (.A(net753),
    .X(net48));
 sky130_fd_sc_hd__buf_1 c710 (.A(net801),
    .X(net681));
 sky130_fd_sc_hd__and2_0 c711 (.A(net1040),
    .B(net677),
    .X(net682));
 sky130_fd_sc_hd__sdfxbp_1 c712 (.CLK(clknet_4_10_0_clk),
    .D(net679),
    .SCD(clknet_1_1__leaf_net678),
    .SCE(net680),
    .Q(net684),
    .Q_N(net683));
 sky130_fd_sc_hd__and3_1 c713 (.A(clknet_1_1__leaf_net678),
    .B(net675),
    .C(net683),
    .X(net685));
 sky130_fd_sc_hd__and2_1 c714 (.A(net680),
    .B(net681),
    .X(net686));
 sky130_fd_sc_hd__buf_1 c715 (.A(net786),
    .X(net687));
 sky130_fd_sc_hd__a2111o_1 c716 (.A1(net677),
    .A2(net686),
    .B1(net687),
    .C1(clknet_1_1__leaf_net674),
    .D1(clknet_1_0__leaf_net897),
    .X(net688));
 sky130_fd_sc_hd__and3_1 c717 (.A(net687),
    .B(net681),
    .C(net686),
    .X(net689));
 sky130_fd_sc_hd__and3_1 c718 (.A(net684),
    .B(clknet_1_1__leaf_net678),
    .C(net677),
    .X(net690));
 sky130_fd_sc_hd__and3_1 c719 (.A(clknet_1_0__leaf_net688),
    .B(clknet_1_0__leaf_net690),
    .C(net679),
    .X(net691));
 sky130_fd_sc_hd__and2_0 c72 (.A(net43),
    .B(net47),
    .X(net49));
 sky130_fd_sc_hd__and3_1 c720 (.A(clknet_1_0__leaf_net690),
    .B(net687),
    .C(net680),
    .X(net692));
 sky130_fd_sc_hd__sdfrtp_1 c721 (.CLK(clknet_4_10_0_clk),
    .D(net687),
    .RESET_B(clknet_1_0__leaf_net690),
    .SCD(net686),
    .SCE(net890),
    .Q(net693));
 sky130_fd_sc_hd__and3_1 c722 (.A(clknet_1_0__leaf_net688),
    .B(net686),
    .C(net693),
    .X(net694));
 sky130_fd_sc_hd__a2111o_1 c723 (.A1(net693),
    .A2(net689),
    .B1(net687),
    .C1(clknet_1_1__leaf_net690),
    .D1(net683),
    .X(net695));
 sky130_fd_sc_hd__mux4_2 c724 (.A0(clknet_1_1__leaf_net694),
    .A1(net693),
    .A2(net675),
    .A3(net680),
    .S0(net890),
    .S1(net906),
    .X(net696));
 sky130_fd_sc_hd__mux4_1 c725 (.A0(net684),
    .A1(clknet_1_1__leaf_net690),
    .A2(clknet_1_1__leaf_net688),
    .A3(net568),
    .S0(clknet_1_0__leaf_net694),
    .X(net697));
 sky130_fd_sc_hd__and2_1 c726 (.A(net597),
    .B(net930),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 c727 (.A(net698),
    .X(net699));
 sky130_fd_sc_hd__buf_1 c728 (.A(net698),
    .X(net700));
 sky130_fd_sc_hd__buf_1 c729 (.A(net699),
    .X(net701));
 sky130_fd_sc_hd__and2_1 c73 (.A(net45),
    .B(net47),
    .X(net50));
 sky130_fd_sc_hd__buf_1 c730 (.A(clknet_1_1__leaf_net961),
    .X(net702));
 sky130_fd_sc_hd__buf_1 c731 (.A(net882),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_1 c732 (.A(net881),
    .X(net704));
 sky130_fd_sc_hd__and2_0 c733 (.A(net700),
    .B(net703),
    .X(net705));
 sky130_fd_sc_hd__and2_0 c734 (.A(net704),
    .B(net703),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 c735 (.A(net771),
    .X(net707));
 sky130_fd_sc_hd__and2_0 c736 (.A(net707),
    .B(net706),
    .X(net708));
 sky130_fd_sc_hd__and2_1 c737 (.A(net682),
    .B(net708),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 c738 (.A(net829),
    .X(net710));
 sky130_fd_sc_hd__buf_1 c739 (.A(net774),
    .X(net711));
 sky130_fd_sc_hd__buf_1 c74 (.A(net1026),
    .X(net51));
 sky130_fd_sc_hd__and2_1 c740 (.A(net710),
    .B(net708),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 c741 (.A(net959),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_1 c742 (.A(net828),
    .X(net714));
 sky130_fd_sc_hd__and2_0 c743 (.A(net713),
    .B(net714),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_1 c744 (.A(net825),
    .X(net716));
 sky130_fd_sc_hd__and3_1 c745 (.A(net715),
    .B(net700),
    .C(net714),
    .X(net717));
 sky130_fd_sc_hd__mux4_1 c746 (.A0(net711),
    .A1(net716),
    .A2(net714),
    .A3(net597),
    .S0(net606),
    .S1(net703),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 c747 (.A(net792),
    .X(net719));
 sky130_fd_sc_hd__buf_1 c748 (.A(clknet_1_1__leaf_net941),
    .X(net720));
 sky130_fd_sc_hd__and2_0 c749 (.A(clknet_1_1__leaf_net720),
    .B(net992),
    .X(net721));
 sky130_fd_sc_hd__dlymetal6s2s_1 c75 (.A(net47),
    .X(net52));
 sky130_fd_sc_hd__and3_1 c750 (.A(net992),
    .B(clknet_1_1__leaf_net721),
    .C(clknet_1_1__leaf_net720),
    .X(net722));
 sky130_fd_sc_hd__or4bb_1 c751 (.A(clknet_1_0__leaf_net721),
    .B(net719),
    .C_N(clknet_1_1__leaf_net722),
    .D_N(net626),
    .X(net723));
 sky130_fd_sc_hd__buf_1 c752 (.A(clknet_1_0__leaf_net941),
    .X(net724));
 sky130_fd_sc_hd__sdfbbn_1 c753 (.CLK_N(clknet_4_10_0_clk),
    .D(clknet_1_1__leaf_net723),
    .RESET_B(clknet_1_1__leaf_net724),
    .SCD(clknet_1_0__leaf_net720),
    .SCE(clknet_1_1__leaf_net722),
    .SET_B(clknet_1_1__leaf_net721),
    .Q(net726),
    .Q_N(net725));
 sky130_fd_sc_hd__a2111o_1 c754 (.A1(net675),
    .A2(clknet_1_1__leaf_net724),
    .B1(clknet_1_0__leaf_net722),
    .C1(net719),
    .D1(net725),
    .X(net727));
 sky130_fd_sc_hd__a2111o_1 c755 (.A1(clknet_1_1__leaf_net727),
    .A2(net726),
    .B1(clknet_1_0__leaf_net723),
    .C1(clknet_1_0__leaf_net724),
    .D1(clknet_1_0__leaf_net722),
    .X(net728));
 sky130_fd_sc_hd__a2111o_1 c756 (.A1(clknet_1_0__leaf_net724),
    .A2(clknet_1_0__leaf_net722),
    .B1(clknet_1_0__leaf_net723),
    .C1(clknet_1_0__leaf_net727),
    .D1(net906),
    .X(net729));
 sky130_fd_sc_hd__buf_1 c76 (.A(net775),
    .X(net53));
 sky130_fd_sc_hd__and3_1 c77 (.A(net49),
    .B(net51),
    .C(net41),
    .X(net54));
 sky130_fd_sc_hd__and2_1 c78 (.A(net53),
    .B(net875),
    .X(net55));
 sky130_fd_sc_hd__and3_1 c79 (.A(net45),
    .B(net55),
    .C(net46),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 c80 (.A(net789),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 c81 (.A(net924),
    .X(net58));
 sky130_fd_sc_hd__and3_1 c82 (.A(net52),
    .B(net53),
    .C(net51),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 c83 (.A(net818),
    .X(net60));
 sky130_fd_sc_hd__and3_1 c84 (.A(net57),
    .B(net56),
    .C(net48),
    .X(net61));
 sky130_fd_sc_hd__buf_1 c85 (.A(net824),
    .X(net62));
 sky130_fd_sc_hd__and3_1 c86 (.A(net48),
    .B(net61),
    .C(net62),
    .X(net63));
 sky130_fd_sc_hd__a2111o_1 c87 (.A1(net46),
    .A2(net62),
    .B1(net51),
    .C1(net56),
    .D1(net923),
    .X(net64));
 sky130_fd_sc_hd__buf_1 c88 (.A(net55),
    .X(net65));
 sky130_fd_sc_hd__and2_0 c89 (.A(net65),
    .B(net1061),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 c90 (.A(net65),
    .X(net67));
 sky130_fd_sc_hd__buf_1 c91 (.A(net56),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 c92 (.A(net919),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 c93 (.A(net919),
    .X(net70));
 sky130_fd_sc_hd__buf_1 c94 (.A(net782),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 c95 (.A(net909),
    .X(net72));
 sky130_fd_sc_hd__and2_1 c96 (.A(net71),
    .B(net1000),
    .X(net73));
 sky130_fd_sc_hd__and2_0 c97 (.A(net70),
    .B(net71),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 c98 (.A(net781),
    .X(net75));
 sky130_fd_sc_hd__and2_0 c99 (.A(net60),
    .B(net71),
    .X(net76));
 sky130_fd_sc_hd__sdfsbp_1 merge757 (.CLK(clknet_4_8_0_clk),
    .D(net646),
    .SCD(net655),
    .SCE(net658),
    .Q(net656),
    .Q_N(net730));
 sky130_fd_sc_hd__buf_1 merge758 (.A(net965),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 merge759 (.A(net850),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 merge760 (.A(net778),
    .X(net734));
 sky130_fd_sc_hd__sdfsbp_1 merge761 (.CLK(clknet_4_0_0_clk),
    .D(net253),
    .SCD(net387),
    .SCE(net386),
    .SET_B(net393),
    .Q(net736),
    .Q_N(net735));
 sky130_fd_sc_hd__clkbuf_1 merge762 (.A(net772),
    .X(net737));
 sky130_fd_sc_hd__buf_1 merge763 (.A(net953),
    .X(net738));
 sky130_fd_sc_hd__or4bb_1 merge764 (.A(clknet_1_0__leaf_net694),
    .B(net606),
    .C_N(clknet_1_0__leaf_net702),
    .D_N(net701),
    .X(net739));
 sky130_fd_sc_hd__sdfxbp_1 merge765 (.CLK(clknet_4_1_0_clk),
    .D(net2),
    .SCD(net985),
    .SCE(net534),
    .Q(net741),
    .Q_N(net740));
 sky130_fd_sc_hd__buf_1 merge766 (.A(net967),
    .X(net742));
 sky130_fd_sc_hd__sdfstp_1 merge767 (.CLK(clknet_4_4_0_clk),
    .D(net22),
    .SCD(net23),
    .SCE(net27),
    .SET_B(net25),
    .Q(net743));
 sky130_fd_sc_hd__sdfstp_1 merge768 (.CLK(clknet_4_14_0_clk),
    .D(net381),
    .SCD(net249),
    .SCE(clknet_1_1__leaf_net501),
    .SET_B(clknet_1_1__leaf_net503),
    .Q(net744));
 sky130_fd_sc_hd__buf_1 merge769 (.A(net1037),
    .X(net745));
 sky130_fd_sc_hd__sdfstp_1 merge770 (.CLK(clknet_4_9_0_clk),
    .D(net564),
    .SCD(net477),
    .SCE(net591),
    .SET_B(net593),
    .Q(net746));
 sky130_fd_sc_hd__sdfxtp_1 merge771 (.CLK(clknet_4_5_0_clk),
    .D(net158),
    .SCD(net159),
    .SCE(net157),
    .Q(net747));
 sky130_fd_sc_hd__clkbuf_1 merge772 (.A(net797),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 merge773 (.A(net951),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 merge774 (.A(net968),
    .X(net750));
 sky130_fd_sc_hd__buf_1 merge775 (.A(clknet_1_1__leaf_net962),
    .X(net751));
 sky130_fd_sc_hd__mux4_1 merge776 (.A0(net717),
    .A1(net626),
    .A2(clknet_1_1__leaf_net722),
    .A3(clknet_1_0__leaf_net720),
    .S0(clknet_1_0__leaf_net721),
    .S1(clknet_1_1__leaf_net723),
    .X(net752));
 sky130_fd_sc_hd__sdfxtp_1 merge777 (.CLK(clknet_4_7_0_clk),
    .D(net44),
    .SCD(net34),
    .SCE(net43),
    .Q(net753));
 sky130_fd_sc_hd__or4bb_1 merge778 (.A(net253),
    .B(net276),
    .C_N(net277),
    .D_N(net928),
    .X(net754));
 sky130_fd_sc_hd__sdfxtp_1 merge779 (.CLK(clknet_4_4_0_clk),
    .D(net296),
    .SCD(net297),
    .SCE(net300),
    .Q(net755));
 sky130_fd_sc_hd__and3_1 merge780 (.A(net42),
    .B(net68),
    .C(net67),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 merge781 (.A(net804),
    .X(net757));
 sky130_fd_sc_hd__dfbbn_1 merge782 (.CLK_N(clknet_4_15_0_clk),
    .D(net226),
    .RESET_B(net89),
    .SET_B(net228),
    .Q(net759),
    .Q_N(net758));
 sky130_fd_sc_hd__buf_1 merge783 (.A(net949),
    .X(net760));
 sky130_fd_sc_hd__sedfxbp_1 merge784 (.CLK(clknet_4_6_0_clk),
    .D(net299),
    .DE(net315),
    .SCD(net64),
    .SCE(net312),
    .Q(net762),
    .Q_N(net761));
 sky130_fd_sc_hd__or4bb_1 merge785 (.A(net116),
    .B(net115),
    .C_N(net114),
    .D_N(net975),
    .X(net763));
 sky130_fd_sc_hd__buf_1 merge786 (.A(net772),
    .X(net764));
 sky130_fd_sc_hd__buf_1 merge787 (.A(net791),
    .X(net765));
 sky130_fd_sc_hd__dfbbn_1 merge788 (.CLK_N(clknet_4_8_0_clk),
    .D(net629),
    .RESET_B(net627),
    .Q(net630),
    .Q_N(net766));
 sky130_fd_sc_hd__dfbbp_1 merge789 (.CLK(clknet_4_11_0_clk),
    .D(net600),
    .RESET_B(net608),
    .SET_B(net994),
    .Q(net769),
    .Q_N(net768));
 sky130_fd_sc_hd__sedfxbp_1 merge790 (.CLK(clknet_4_11_0_clk),
    .D(net701),
    .DE(clknet_1_1__leaf_net702),
    .SCD(net619),
    .SCE(net613),
    .Q(net771),
    .Q_N(net770));
 sky130_fd_sc_hd__sedfxtp_2 merge791 (.CLK(clknet_4_12_0_clk),
    .D(net180),
    .DE(net181),
    .SCD(net134),
    .SCE(net136),
    .Q(net772));
 sky130_fd_sc_hd__sedfxtp_1 merge792 (.CLK(clknet_4_0_0_clk),
    .D(net261),
    .DE(net258),
    .SCD(net118),
    .SCE(net116),
    .Q(net773));
 sky130_fd_sc_hd__sedfxtp_1 merge793 (.CLK(clknet_4_8_0_clk),
    .D(net709),
    .DE(net700),
    .SCD(net570),
    .SCE(net576),
    .Q(net774));
 sky130_fd_sc_hd__sdfrbp_1 merge794 (.CLK(clknet_4_7_0_clk),
    .D(net79),
    .RESET_B(net47),
    .SCD(net49),
    .SCE(clknet_1_0__leaf_net895),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__sdfrbp_1 merge795 (.CLK(clknet_4_1_0_clk),
    .D(net253),
    .RESET_B(net1003),
    .SCD(net298),
    .SCE(net300),
    .Q(net778),
    .Q_N(net777));
 sky130_fd_sc_hd__sdfrtn_1 merge796 (.CLK_N(clknet_4_9_0_clk),
    .D(net433),
    .RESET_B(net1044),
    .SCD(net476),
    .SCE(net475),
    .Q(net779));
 sky130_fd_sc_hd__or4bb_1 merge797 (.A(net344),
    .B(net345),
    .C_N(net66),
    .D_N(net68),
    .X(net780));
 sky130_fd_sc_hd__sdfxbp_1 merge798 (.CLK(clknet_4_7_0_clk),
    .D(net65),
    .SCD(net68),
    .SCE(net73),
    .Q(net782),
    .Q_N(net781));
 sky130_fd_sc_hd__sdfrtp_1 merge799 (.CLK(clknet_4_7_0_clk),
    .D(net50),
    .RESET_B(net44),
    .SCD(net26),
    .SCE(net27),
    .Q(net783));
 sky130_fd_sc_hd__or4bb_1 merge800 (.A(net115),
    .B(net116),
    .C_N(net138),
    .D_N(net136),
    .X(net784));
 sky130_fd_sc_hd__or4bb_1 merge801 (.A(net279),
    .B(net286),
    .C_N(net51),
    .D_N(net52),
    .X(net785));
 sky130_fd_sc_hd__sdfrtp_1 merge802 (.CLK(clknet_4_9_0_clk),
    .D(net416),
    .RESET_B(net419),
    .SCD(net685),
    .SCE(clknet_1_0__leaf_net678),
    .Q(net786));
 sky130_fd_sc_hd__sdfrtp_1 merge803 (.CLK(clknet_4_11_0_clk),
    .D(net607),
    .RESET_B(net1014),
    .SCD(net499),
    .SCE(net997),
    .Q(net787));
 sky130_fd_sc_hd__or4bb_1 merge804 (.A(net119),
    .B(clknet_1_0__leaf_net142),
    .C_N(net135),
    .D_N(net880),
    .X(net788));
 sky130_fd_sc_hd__sdfsbp_1 merge805 (.CLK(clknet_4_7_0_clk),
    .D(net75),
    .SCD(net79),
    .SCE(net53),
    .SET_B(net52),
    .Q(net790),
    .Q_N(net789));
 sky130_fd_sc_hd__buf_1 merge806 (.A(net958),
    .X(net791));
 sky130_fd_sc_hd__sdfsbp_1 merge807 (.CLK(clknet_4_9_0_clk),
    .D(net439),
    .SCD(net438),
    .SCE(net705),
    .SET_B(net1001),
    .Q(net793),
    .Q_N(net792));
 sky130_fd_sc_hd__buf_1 merge808 (.A(net957),
    .X(net794));
 sky130_fd_sc_hd__sdfstp_1 merge809 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net503),
    .SCD(clknet_1_0__leaf_net501),
    .SCE(net994),
    .SET_B(net484),
    .Q(net795));
 sky130_fd_sc_hd__sdfstp_1 merge810 (.CLK(clknet_4_2_0_clk),
    .D(net544),
    .SCD(net541),
    .SCE(net513),
    .SET_B(net519),
    .Q(net796));
 sky130_fd_sc_hd__sdfstp_1 merge811 (.CLK(clknet_4_7_0_clk),
    .D(net201),
    .SCD(net202),
    .SCE(net166),
    .SET_B(net160),
    .Q(net797));
 sky130_fd_sc_hd__sedfxbp_1 merge812 (.CLK(clknet_4_2_0_clk),
    .D(net519),
    .DE(net516),
    .SCD(net1033),
    .SCE(net521),
    .Q(net799),
    .Q_N(net798));
 sky130_fd_sc_hd__sedfxbp_1 merge813 (.CLK(clknet_4_10_0_clk),
    .D(net568),
    .DE(net680),
    .SCD(net441),
    .SCE(net438),
    .Q(net801),
    .Q_N(net800));
 sky130_fd_sc_hd__sedfxtp_1 merge814 (.CLK(clknet_4_2_0_clk),
    .D(net254),
    .DE(net251),
    .SCD(net541),
    .SCE(net885),
    .Q(net802));
 sky130_fd_sc_hd__sedfxtp_2 merge815 (.CLK(clknet_4_14_0_clk),
    .D(net357),
    .DE(net504),
    .SCD(clknet_1_1__leaf_net503),
    .SCE(clknet_1_1__leaf_net932),
    .Q(net803));
 sky130_fd_sc_hd__sedfxtp_1 merge816 (.CLK(clknet_4_3_0_clk),
    .D(net254),
    .DE(net410),
    .SCD(net416),
    .SCE(net929),
    .Q(net804));
 sky130_fd_sc_hd__sdfrbp_1 merge817 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_0__leaf_net370),
    .RESET_B(clknet_1_0__leaf_net366),
    .SCD(net480),
    .SCE(net994),
    .Q(net806),
    .Q_N(net805));
 sky130_fd_sc_hd__sdfrbp_1 merge818 (.CLK(clknet_4_8_0_clk),
    .D(net660),
    .RESET_B(net657),
    .SCD(net545),
    .SCE(net541),
    .Q(net808),
    .Q_N(net807));
 sky130_fd_sc_hd__sdfrtn_1 merge819 (.CLK_N(clknet_4_8_0_clk),
    .D(net410),
    .RESET_B(net514),
    .SCD(net664),
    .SCE(net665),
    .Q(net809));
 sky130_fd_sc_hd__sdfrtp_1 merge820 (.CLK(clknet_4_9_0_clk),
    .D(net438),
    .RESET_B(net1006),
    .SCD(net479),
    .SCE(net489),
    .Q(net810));
 sky130_fd_sc_hd__sdfrtp_1 merge821 (.CLK(clknet_4_6_0_clk),
    .D(net413),
    .RESET_B(net410),
    .SCD(net459),
    .SCE(net470),
    .Q(net811));
 sky130_fd_sc_hd__sdfrtp_1 merge822 (.CLK(clknet_4_3_0_clk),
    .D(net277),
    .RESET_B(net291),
    .SCD(net447),
    .SCE(net446),
    .Q(net812));
 sky130_fd_sc_hd__sdfsbp_1 merge823 (.CLK(clknet_4_5_0_clk),
    .D(net172),
    .SCE(net159),
    .SET_B(net888),
    .Q(net173),
    .Q_N(net813));
 sky130_fd_sc_hd__or4bb_1 merge824 (.A(net493),
    .B(net321),
    .C_N(net323),
    .X(net815));
 sky130_fd_sc_hd__sdfsbp_1 merge825 (.CLK(clknet_4_12_0_clk),
    .D(net322),
    .SCD(net318),
    .SCE(net489),
    .SET_B(net490),
    .Q(net817),
    .Q_N(net816));
 sky130_fd_sc_hd__sdfstp_1 merge826 (.CLK(clknet_4_6_0_clk),
    .D(net58),
    .SCD(net50),
    .SCE(net460),
    .SET_B(net1055),
    .Q(net818));
 sky130_fd_sc_hd__sdfstp_1 merge827 (.CLK(clknet_4_12_0_clk),
    .D(net327),
    .SCD(net330),
    .SCE(net371),
    .SET_B(clknet_1_0__leaf_net370),
    .Q(net819));
 sky130_fd_sc_hd__sdfstp_1 merge828 (.CLK(clknet_4_10_0_clk),
    .D(net653),
    .SCD(net662),
    .SCE(net632),
    .SET_B(net629),
    .Q(net820));
 sky130_fd_sc_hd__sedfxbp_1 merge829 (.CLK(clknet_4_8_0_clk),
    .D(net661),
    .DE(net658),
    .SCD(net487),
    .SCE(net994),
    .Q(net822),
    .Q_N(net821));
 sky130_fd_sc_hd__sedfxbp_1 merge830 (.CLK(clknet_4_7_0_clk),
    .D(net50),
    .DE(net48),
    .SCD(net202),
    .SCE(net207),
    .Q(net824),
    .Q_N(net823));
 sky130_fd_sc_hd__sedfxtp_1 merge831 (.CLK(clknet_4_10_0_clk),
    .D(net633),
    .DE(net629),
    .SCD(net706),
    .SCE(net606),
    .Q(net825));
 sky130_fd_sc_hd__sedfxtp_1 merge832 (.CLK(clknet_4_14_0_clk),
    .D(clknet_1_1__leaf_net370),
    .DE(clknet_1_0__leaf_net374),
    .SCD(net182),
    .SCE(net186),
    .Q(net826));
 sky130_fd_sc_hd__sedfxtp_1 merge833 (.CLK(clknet_4_14_0_clk),
    .D(net182),
    .DE(net184),
    .SCD(net367),
    .SCE(clknet_1_0__leaf_net368),
    .Q(net827));
 sky130_fd_sc_hd__sdfrbp_1 merge834 (.CLK(clknet_4_8_0_clk),
    .D(net703),
    .RESET_B(net1041),
    .SCD(net698),
    .SCE(net701),
    .Q(net829),
    .Q_N(net828));
 sky130_fd_sc_hd__mux4_1 merge835 (.A0(net114),
    .A1(net119),
    .A2(net113),
    .A3(clknet_1_0__leaf_net121),
    .S0(net124),
    .S1(net116),
    .X(net830));
 sky130_fd_sc_hd__sdfrbp_1 merge836 (.CLK(clknet_4_13_0_clk),
    .D(net185),
    .RESET_B(net187),
    .SCD(net91),
    .SCE(net88),
    .Q(net832),
    .Q_N(net831));
 sky130_fd_sc_hd__mux4_1 merge837 (.A0(net451),
    .A1(net450),
    .A2(net446),
    .A3(net665),
    .S0(net671),
    .S1(clknet_1_0__leaf_net940),
    .X(net833));
 sky130_fd_sc_hd__mux4_1 merge838 (.A0(net457),
    .A1(net462),
    .A2(net464),
    .A3(net482),
    .S0(net489),
    .S1(net490),
    .X(net834));
 sky130_fd_sc_hd__mux4_1 merge839 (.A0(net300),
    .A1(net252),
    .A2(net254),
    .A3(net251),
    .S0(net867),
    .S1(net937),
    .X(net835));
 sky130_fd_sc_hd__mux4_1 merge840 (.A0(net297),
    .A1(net300),
    .A2(net302),
    .A3(net460),
    .S0(net458),
    .S1(net321),
    .X(net836));
 sky130_fd_sc_hd__mux4_1 merge841 (.A0(net125),
    .A1(clknet_1_1__leaf_net121),
    .A2(net116),
    .A3(net258),
    .S0(net259),
    .S1(net253),
    .X(net837));
 sky130_fd_sc_hd__mux4_1 merge842 (.A0(net662),
    .A1(clknet_1_0__leaf_net678),
    .A2(net500),
    .A3(clknet_1_0__leaf_net365),
    .S0(clknet_1_0__leaf_net503),
    .S1(clknet_1_1__leaf_net897),
    .X(net838));
 sky130_fd_sc_hd__mux4_1 merge843 (.A0(net273),
    .A1(net289),
    .A2(net278),
    .A3(net333),
    .S0(net328),
    .S1(net299),
    .X(net839));
 sky130_fd_sc_hd__mux4_1 merge844 (.A0(net535),
    .A1(net541),
    .A2(net543),
    .A3(net30),
    .S0(net20),
    .S1(net27),
    .X(net840));
 sky130_fd_sc_hd__mux4_1 merge845 (.A0(net585),
    .A1(net587),
    .A2(net590),
    .A3(net257),
    .S0(net265),
    .S1(net263),
    .X(net841));
 sky130_fd_sc_hd__sdfrtn_1 merge846 (.CLK_N(clknet_4_13_0_clk),
    .D(net236),
    .RESET_B(net1007),
    .SCD(net98),
    .SCE(net72),
    .Q(net842));
 sky130_fd_sc_hd__mux4_1 merge847 (.A0(net458),
    .A1(net460),
    .A2(net464),
    .A3(net511),
    .S0(clknet_1_1__leaf_net503),
    .S1(net901),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 merge848 (.A0(net167),
    .A1(net172),
    .A2(net173),
    .A3(net479),
    .S0(net207),
    .S1(net206),
    .X(net844));
 sky130_fd_sc_hd__or4bb_1 merge849 (.A(net226),
    .B(net228),
    .C_N(net100),
    .D_N(net98),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 merge850 (.A0(net281),
    .A1(net283),
    .A2(net273),
    .A3(net577),
    .S0(net578),
    .S1(clknet_1_0__leaf_net579),
    .X(net846));
 sky130_fd_sc_hd__mux4_1 merge851 (.A0(net544),
    .A1(net551),
    .A2(net542),
    .A3(net712),
    .S0(net709),
    .S1(net711),
    .X(net847));
 sky130_fd_sc_hd__mux4_1 merge852 (.A0(net462),
    .A1(net464),
    .A2(net470),
    .A3(net505),
    .S0(net996),
    .S1(clknet_1_0__leaf_net503),
    .X(net848));
 sky130_fd_sc_hd__sdfbbn_1 merge853 (.CLK_N(clknet_4_12_0_clk),
    .D(net92),
    .RESET_B(net90),
    .SCD(net468),
    .SCE(net464),
    .SET_B(net470),
    .Q(net850),
    .Q_N(net849));
 sky130_fd_sc_hd__mux4_1 merge854 (.A0(net673),
    .A1(net671),
    .A2(net699),
    .A3(net597),
    .S0(net606),
    .S1(clknet_1_1__leaf_net940),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 merge855 (.A0(net189),
    .A1(net180),
    .A2(net191),
    .A3(clknet_1_0__leaf_net368),
    .S0(net363),
    .S1(net346),
    .X(net852));
 sky130_fd_sc_hd__sdfbbp_1 merge856 (.CLK(clknet_4_4_0_clk),
    .D(net25),
    .RESET_B(net27),
    .SCD(net983),
    .SCE(net32),
    .SET_B(net30),
    .Q(net854),
    .Q_N(net853));
 sky130_fd_sc_hd__mux4_1 merge857 (.A0(net571),
    .A1(net575),
    .A2(net572),
    .A3(net981),
    .S0(net139),
    .S1(net136),
    .X(net855));
 sky130_fd_sc_hd__mux4_1 merge858 (.A0(net431),
    .A1(net435),
    .A2(net436),
    .A3(net390),
    .S0(net395),
    .S1(net394),
    .X(net856));
 sky130_fd_sc_hd__mux4_1 merge859 (.A0(net557),
    .A1(net568),
    .A2(net556),
    .A3(net491),
    .S0(clknet_1_0__leaf_net503),
    .S1(clknet_1_0__leaf_net365),
    .X(net857));
 sky130_fd_sc_hd__mux4_1 merge860 (.A0(net29),
    .A1(net31),
    .A2(net32),
    .A3(net343),
    .S0(net330),
    .S1(net339),
    .X(net858));
 sky130_fd_sc_hd__mux4_1 merge861 (.A0(net419),
    .A1(net425),
    .A2(net426),
    .A3(net263),
    .S0(net265),
    .S1(net929),
    .X(net859));
 sky130_fd_sc_hd__dfrbp_1 merge862 (.CLK(clknet_4_15_0_clk),
    .D(net240),
    .RESET_B(net247),
    .Q(net861),
    .Q_N(net860));
 sky130_fd_sc_hd__and2_0 merge863 (.A(net729),
    .B(net728),
    .X(net862));
 sky130_fd_sc_hd__dfrbp_1 merge864 (.CLK(clknet_4_0_0_clk),
    .D(net270),
    .Q(net271),
    .Q_N(net863));
 sky130_fd_sc_hd__and2_0 merge865 (.A(net355),
    .B(net362),
    .X(net865));
 sky130_fd_sc_hd__dfrtn_1 merge866 (.CLK_N(clknet_4_15_0_clk),
    .D(net372),
    .RESET_B(net383),
    .Q(net866));
 sky130_fd_sc_hd__dfrtp_1 merge867 (.CLK(clknet_4_1_0_clk),
    .D(net304),
    .RESET_B(net310),
    .Q(net867));
 sky130_fd_sc_hd__dfrtp_1 merge868 (.CLK(clknet_4_1_0_clk),
    .D(net7),
    .RESET_B(net8),
    .Q(net868));
 sky130_fd_sc_hd__dfrtp_1 merge869 (.CLK(clknet_4_2_0_clk),
    .D(net429),
    .RESET_B(net432),
    .Q(net869));
 sky130_fd_sc_hd__dfsbp_1 merge870 (.CLK(clknet_4_5_0_clk),
    .D(net38),
    .SET_B(net1049),
    .Q(net871),
    .Q_N(net870));
 sky130_fd_sc_hd__dfsbp_1 merge871 (.CLK(clknet_4_11_0_clk),
    .D(net622),
    .SET_B(net623),
    .Q(net873),
    .Q_N(net872));
 sky130_fd_sc_hd__dfstp_1 merge872 (.CLK(clknet_4_8_0_clk),
    .D(net645),
    .SET_B(net652),
    .Q(net874));
 sky130_fd_sc_hd__dfstp_1 merge873 (.CLK(clknet_4_7_0_clk),
    .D(net54),
    .SET_B(net59),
    .Q(net875));
 sky130_fd_sc_hd__dfstp_1 merge874 (.CLK(clknet_4_9_0_clk),
    .D(net448),
    .SET_B(net454),
    .Q(net876));
 sky130_fd_sc_hd__dlrbn_1 merge875 (.D(net143),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net154),
    .Q(net878),
    .Q_N(net877));
 sky130_fd_sc_hd__dlrbn_1 merge876 (.D(net127),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net763),
    .Q(net880),
    .Q_N(net879));
 sky130_fd_sc_hd__dlrbp_1 merge877 (.D(net718),
    .GATE(clknet_4_9_0_clk),
    .RESET_B(net739),
    .Q(net882),
    .Q_N(net881));
 sky130_fd_sc_hd__dlrbp_1 merge878 (.D(net214),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net217),
    .Q(net884),
    .Q_N(net883));
 sky130_fd_sc_hd__dlrtn_1 merge879 (.D(net549),
    .GATE_N(clknet_4_2_0_clk),
    .RESET_B(net555),
    .Q(net885));
 sky130_fd_sc_hd__and2_0 merge880 (.A(net495),
    .B(net496),
    .X(net886));
 sky130_fd_sc_hd__dlrtn_1 merge881 (.D(net197),
    .GATE_N(clknet_4_15_0_clk),
    .Q(net198));
 sky130_fd_sc_hd__dlrtn_1 merge882 (.GATE_N(clknet_4_5_0_clk),
    .RESET_B(net169),
    .Q(net170));
 sky130_fd_sc_hd__dlrtp_1 merge883 (.D(net404),
    .GATE(clknet_4_2_0_clk),
    .RESET_B(net407),
    .Q(net889));
 sky130_fd_sc_hd__dlrtp_1 merge884 (.D(net691),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net692),
    .Q(net890));
 sky130_fd_sc_hd__dlrtp_1 merge885 (.D(net666),
    .GATE(clknet_4_8_0_clk),
    .RESET_B(net669),
    .Q(net891));
 sky130_fd_sc_hd__edfxbp_1 merge886 (.CLK(clknet_4_3_0_clk),
    .D(net290),
    .DE(net294),
    .Q(net893),
    .Q_N(net892));
 sky130_fd_sc_hd__edfxtp_1 merge887 (.CLK(clknet_4_12_0_clk),
    .D(net324),
    .DE(net334),
    .Q(net894));
 sky130_fd_sc_hd__sdlclkp_1 merge888 (.CLK(clknet_4_13_0_clk),
    .GATE(net80),
    .SCE(net82),
    .GCLK(net895));
 sky130_fd_sc_hd__sdlclkp_2 merge889 (.CLK(clknet_4_11_0_clk),
    .GATE(net473),
    .SCE(net478),
    .GCLK(net998));
 sky130_fd_sc_hd__and2_0 merge890 (.A(net530),
    .B(net533),
    .X(net896));
 sky130_fd_sc_hd__sdlclkp_4 merge891 (.CLK(clknet_4_9_0_clk),
    .GATE(net581),
    .GCLK(net897));
 sky130_fd_sc_hd__and2_0 merge892 (.A(net108),
    .B(net109),
    .X(net898));
 sky130_fd_sc_hd__dfrbp_1 merge893 (.CLK(clknet_4_9_0_clk),
    .D(net594),
    .RESET_B(net1023),
    .Q(net900),
    .Q_N(net899));
 sky130_fd_sc_hd__dfrbp_1 merge894 (.CLK(clknet_4_14_0_clk),
    .D(net507),
    .RESET_B(net509),
    .Q(net902),
    .Q_N(net901));
 sky130_fd_sc_hd__dfrtn_1 merge895 (.CLK_N(clknet_4_3_0_clk),
    .D(net408),
    .RESET_B(net155),
    .Q(net903));
 sky130_fd_sc_hd__dfrtp_1 merge896 (.CLK(clknet_4_4_0_clk),
    .D(net14),
    .RESET_B(net16),
    .Q(net904));
 sky130_fd_sc_hd__dfrtp_1 merge897 (.CLK(clknet_4_2_0_clk),
    .D(net409),
    .RESET_B(net560),
    .Q(net905));
 sky130_fd_sc_hd__dfrtp_1 merge898 (.CLK(clknet_4_10_0_clk),
    .D(net695),
    .RESET_B(net862),
    .Q(net906));
 sky130_fd_sc_hd__dfsbp_1 merge899 (.CLK(clknet_4_11_0_clk),
    .D(net618),
    .Q(net624),
    .Q_N(net907));
 sky130_fd_sc_hd__dfsbp_1 merge900 (.CLK(clknet_4_6_0_clk),
    .D(net338),
    .SET_B(net780),
    .Q(net910),
    .Q_N(net909));
 sky130_fd_sc_hd__dfstp_1 merge901 (.CLK(clknet_4_15_0_clk),
    .D(net220),
    .SET_B(net385),
    .Q(net911));
 sky130_fd_sc_hd__dfstp_1 merge902 (.CLK(clknet_4_13_0_clk),
    .D(net19),
    .SET_B(net199),
    .Q(net912));
 sky130_fd_sc_hd__dfstp_1 merge903 (.CLK(clknet_4_15_0_clk),
    .D(net221),
    .SET_B(net384),
    .Q(net913));
 sky130_fd_sc_hd__dlrbn_1 merge904 (.D(net224),
    .GATE_N(clknet_4_5_0_clk),
    .RESET_B(net1036),
    .Q(net915),
    .Q_N(net914));
 sky130_fd_sc_hd__dlrbn_1 merge905 (.D(net845),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net219),
    .Q(net917),
    .Q_N(net916));
 sky130_fd_sc_hd__dlrbp_1 merge906 (.D(net756),
    .GATE(clknet_4_13_0_clk),
    .RESET_B(net898),
    .Q(net919),
    .Q_N(net918));
 sky130_fd_sc_hd__dlrbp_1 merge907 (.D(net149),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net156),
    .Q(net921),
    .Q_N(net920));
 sky130_fd_sc_hd__dlrtn_1 merge908 (.D(net754),
    .GATE_N(clknet_4_3_0_clk),
    .RESET_B(net846),
    .Q(net922));
 sky130_fd_sc_hd__dlrtn_1 merge909 (.D(net63),
    .GATE_N(clknet_4_13_0_clk),
    .RESET_B(net865),
    .Q(net923));
 sky130_fd_sc_hd__dlrtn_1 merge910 (.D(net285),
    .GATE_N(clknet_4_6_0_clk),
    .RESET_B(net785),
    .Q(net924));
 sky130_fd_sc_hd__dlrtp_1 merge911 (.D(net4),
    .GATE(clknet_4_1_0_clk),
    .RESET_B(net17),
    .Q(net925));
 sky130_fd_sc_hd__dlrtp_1 merge912 (.GATE(clknet_4_14_0_clk),
    .RESET_B(net886),
    .Q(net815));
 sky130_fd_sc_hd__dlrtp_1 merge913 (.GATE(clknet_4_8_0_clk),
    .RESET_B(net896),
    .Q(net927));
 sky130_fd_sc_hd__edfxbp_1 merge914 (.CLK(clknet_4_1_0_clk),
    .D(net264),
    .DE(net272),
    .Q(net929),
    .Q_N(net928));
 sky130_fd_sc_hd__edfxtp_1 merge915 (.CLK(clknet_4_10_0_clk),
    .D(net696),
    .Q(net697));
 sky130_fd_sc_hd__sdlclkp_1 merge916 (.CLK(clknet_4_1_0_clk),
    .GATE(net784),
    .SCE(net788),
    .GCLK(net931));
 sky130_fd_sc_hd__sdlclkp_2 merge917 (.CLK(clknet_4_12_0_clk),
    .GATE(net351),
    .SCE(net354),
    .GCLK(net932));
 sky130_fd_sc_hd__dfxbp_1 s918 (.CLK(clknet_4_0_0_clk),
    .D(net132),
    .Q(net934),
    .Q_N(net933));
 sky130_fd_sc_hd__dfxbp_1 s919 (.CLK(clknet_4_1_0_clk),
    .D(net133),
    .Q(net936),
    .Q_N(net935));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_4_0_clk),
    .D(net306),
    .Q(net937));
 sky130_fd_sc_hd__dfxtp_1 s921 (.CLK(clknet_4_6_0_clk),
    .D(net316),
    .Q(net938));
 sky130_fd_sc_hd__dfxtp_1 s922 (.CLK(clknet_4_11_0_clk),
    .D(net598),
    .Q(net939));
 sky130_fd_sc_hd__dlclkp_1 s923 (.CLK(clknet_4_8_0_clk),
    .GATE(net672),
    .GCLK(net940));
 sky130_fd_sc_hd__dlclkp_2 s924 (.CLK(clknet_4_11_0_clk),
    .GATE(net752),
    .GCLK(net941));
 sky130_fd_sc_hd__dlclkp_4 s925 (.CLK(clknet_4_0_0_clk),
    .GATE(net830),
    .GCLK(net942));
 sky130_fd_sc_hd__dlxbn_2 s926 (.D(net833),
    .GATE_N(clknet_4_8_0_clk),
    .Q(net944),
    .Q_N(net943));
 sky130_fd_sc_hd__dlxbn_1 s927 (.D(net834),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net946),
    .Q_N(net945));
 sky130_fd_sc_hd__dlxbp_1 s928 (.D(net835),
    .GATE(clknet_4_3_0_clk),
    .Q(net948),
    .Q_N(net947));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net836),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net949));
 sky130_fd_sc_hd__dlxtn_1 s930 (.D(net837),
    .GATE_N(clknet_4_0_0_clk),
    .Q(net950));
 sky130_fd_sc_hd__dlxtn_1 s931 (.D(net838),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net951));
 sky130_fd_sc_hd__dlxtp_1 s932 (.D(net839),
    .GATE(clknet_4_6_0_clk),
    .Q(net952));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s933 (.D(net840),
    .SLEEP_B(clknet_4_6_0_clk),
    .Q(net953));
 sky130_fd_sc_hd__dfxbp_1 s934 (.CLK(clknet_4_9_0_clk),
    .D(net841),
    .Q(net955),
    .Q_N(net954));
 sky130_fd_sc_hd__dfxbp_1 s935 (.CLK(clknet_4_14_0_clk),
    .D(net843),
    .Q(net957),
    .Q_N(net956));
 sky130_fd_sc_hd__dfxtp_1 s936 (.CLK(clknet_4_7_0_clk),
    .D(net844),
    .Q(net958));
 sky130_fd_sc_hd__dfxtp_1 s937 (.CLK(clknet_4_8_0_clk),
    .D(net847),
    .Q(net959));
 sky130_fd_sc_hd__dfxtp_1 s938 (.CLK(clknet_4_14_0_clk),
    .D(net848),
    .Q(net960));
 sky130_fd_sc_hd__dlclkp_1 s939 (.CLK(clknet_4_10_0_clk),
    .GATE(net851),
    .GCLK(net961));
 sky130_fd_sc_hd__dlclkp_2 s940 (.CLK(clknet_4_15_0_clk),
    .GATE(net852),
    .GCLK(net962));
 sky130_fd_sc_hd__dlclkp_4 s941 (.CLK(clknet_4_3_0_clk),
    .GATE(net855),
    .GCLK(net963));
 sky130_fd_sc_hd__dlxbn_1 s942 (.D(net856),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net965),
    .Q_N(net964));
 sky130_fd_sc_hd__dlxbn_1 s943 (.D(net857),
    .GATE_N(clknet_4_11_0_clk),
    .Q(net967),
    .Q_N(net966));
 sky130_fd_sc_hd__dlxbp_1 s944 (.D(net858),
    .GATE(clknet_4_6_0_clk),
    .Q(net969),
    .Q_N(net968));
 sky130_fd_sc_hd__dlxtn_1 s945 (.D(net859),
    .GATE_N(clknet_4_3_0_clk),
    .Q(net970));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(in1),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in12),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(in17),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(in18),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in21),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in22),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(in23),
    .X(net980));
 sky130_fd_sc_hd__buf_1 input17 (.A(in24),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(in3),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in4),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in5),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(in6),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in7),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in8),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in9),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(clknet_1_1__leaf_net989),
    .X(out11));
 sky130_fd_sc_hd__buf_2 output26 (.A(net990),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output27 (.A(net991),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output28 (.A(net992),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output29 (.A(net993),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output30 (.A(net994),
    .X(out23));
 sky130_fd_sc_hd__clkbuf_4 output31 (.A(net995),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output32 (.A(net996),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output33 (.A(net997),
    .X(out5));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(clknet_1_1__leaf_net998),
    .X(out7));
 sky130_fd_sc_hd__buf_4 output35 (.A(net999),
    .X(out9));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net72),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net963 (.A(net963),
    .X(clknet_0_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_0__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net963 (.A(clknet_0_net963),
    .X(clknet_1_1__leaf_net963));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net579 (.A(net579),
    .X(clknet_0_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_0__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net579 (.A(clknet_0_net579),
    .X(clknet_1_1__leaf_net579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net897 (.A(net897),
    .X(clknet_0_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_0__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net897 (.A(clknet_0_net897),
    .X(clknet_1_1__leaf_net897));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net688 (.A(net688),
    .X(clknet_0_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net688 (.A(clknet_0_net688),
    .X(clknet_1_0__leaf_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net688 (.A(clknet_0_net688),
    .X(clknet_1_1__leaf_net688));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net694 (.A(net694),
    .X(clknet_0_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_0__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net694 (.A(clknet_0_net694),
    .X(clknet_1_1__leaf_net694));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net146 (.A(net146),
    .X(clknet_0_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_0__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net146 (.A(clknet_0_net146),
    .X(clknet_1_1__leaf_net146));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net962 (.A(net962),
    .X(clknet_0_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net962 (.A(clknet_0_net962),
    .X(clknet_1_0__leaf_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net962 (.A(clknet_0_net962),
    .X(clknet_1_1__leaf_net962));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net751 (.A(net751),
    .X(clknet_0_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_0__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net751 (.A(clknet_0_net751),
    .X(clknet_1_1__leaf_net751));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net369 (.A(net369),
    .X(clknet_0_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_0__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net369 (.A(clknet_0_net369),
    .X(clknet_1_1__leaf_net369));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net380 (.A(net380),
    .X(clknet_0_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_0__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net380 (.A(clknet_0_net380),
    .X(clknet_1_1__leaf_net380));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net503 (.A(net503),
    .X(clknet_0_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net503 (.A(clknet_0_net503),
    .X(clknet_1_1__leaf_net503));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net382 (.A(net382),
    .X(clknet_0_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_0__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net382 (.A(clknet_0_net382),
    .X(clknet_1_1__leaf_net382));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net370 (.A(net370),
    .X(clknet_0_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_0__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net370 (.A(clknet_0_net370),
    .X(clknet_1_1__leaf_net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net365 (.A(net365),
    .X(clknet_0_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net365 (.A(clknet_0_net365),
    .X(clknet_1_1__leaf_net365));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net501 (.A(net501),
    .X(clknet_0_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_0__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net501 (.A(clknet_0_net501),
    .X(clknet_1_1__leaf_net501));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net989 (.A(net989),
    .X(clknet_0_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net989 (.A(clknet_0_net989),
    .X(clknet_1_0__leaf_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net989 (.A(clknet_0_net989),
    .X(clknet_1_1__leaf_net989));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net374 (.A(net374),
    .X(clknet_0_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_0__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net374 (.A(clknet_0_net374),
    .X(clknet_1_1__leaf_net374));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net193 (.A(net193),
    .X(clknet_0_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_0__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net193 (.A(clknet_0_net193),
    .X(clknet_1_1__leaf_net193));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net961 (.A(net961),
    .X(clknet_0_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_0__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net961 (.A(clknet_0_net961),
    .X(clknet_1_1__leaf_net961));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net702 (.A(net702),
    .X(clknet_0_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_0__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net702 (.A(clknet_0_net702),
    .X(clknet_1_1__leaf_net702));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net674 (.A(net674),
    .X(clknet_0_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_0__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net674 (.A(clknet_0_net674),
    .X(clknet_1_1__leaf_net674));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net678 (.A(net678),
    .X(clknet_0_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_0__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net678 (.A(clknet_0_net678),
    .X(clknet_1_1__leaf_net678));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net690 (.A(net690),
    .X(clknet_0_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_0__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net690 (.A(clknet_0_net690),
    .X(clknet_1_1__leaf_net690));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net942 (.A(net942),
    .X(clknet_0_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_0__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net942 (.A(clknet_0_net942),
    .X(clknet_1_1__leaf_net942));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net123 (.A(net123),
    .X(clknet_0_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net123 (.A(clknet_0_net123),
    .X(clknet_1_0__leaf_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net123 (.A(clknet_0_net123),
    .X(clknet_1_1__leaf_net123));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net129 (.A(net129),
    .X(clknet_0_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_0__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net129 (.A(clknet_0_net129),
    .X(clknet_1_1__leaf_net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net131 (.A(net131),
    .X(clknet_0_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_0__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net131 (.A(clknet_0_net131),
    .X(clknet_1_1__leaf_net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net941 (.A(net941),
    .X(clknet_0_net941));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net941 (.A(clknet_0_net941),
    .X(clknet_1_0__leaf_net941));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net941 (.A(clknet_0_net941),
    .X(clknet_1_1__leaf_net941));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net724 (.A(net724),
    .X(clknet_0_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_0__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net724 (.A(clknet_0_net724),
    .X(clknet_1_1__leaf_net724));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net727 (.A(net727),
    .X(clknet_0_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_0__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net727 (.A(clknet_0_net727),
    .X(clknet_1_1__leaf_net727));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net720 (.A(net720),
    .X(clknet_0_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_0__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net720 (.A(clknet_0_net720),
    .X(clknet_1_1__leaf_net720));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net722 (.A(net722),
    .X(clknet_0_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net722 (.A(clknet_0_net722),
    .X(clknet_1_0__leaf_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net722 (.A(clknet_0_net722),
    .X(clknet_1_1__leaf_net722));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net723 (.A(net723),
    .X(clknet_0_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net723 (.A(clknet_0_net723),
    .X(clknet_1_0__leaf_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net723 (.A(clknet_0_net723),
    .X(clknet_1_1__leaf_net723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net721 (.A(net721),
    .X(clknet_0_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_0__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net721 (.A(clknet_0_net721),
    .X(clknet_1_1__leaf_net721));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net940 (.A(net940),
    .X(clknet_0_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net940 (.A(clknet_0_net940),
    .X(clknet_1_0__leaf_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net940 (.A(clknet_0_net940),
    .X(clknet_1_1__leaf_net940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net932 (.A(net932),
    .X(clknet_0_net932));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net932 (.A(clknet_0_net932),
    .X(clknet_1_0__leaf_net932));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net932 (.A(clknet_0_net932),
    .X(clknet_1_1__leaf_net932));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net366 (.A(net366),
    .X(clknet_0_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_0__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net366 (.A(clknet_0_net366),
    .X(clknet_1_1__leaf_net366));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net368 (.A(net368),
    .X(clknet_0_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_0__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net368 (.A(clknet_0_net368),
    .X(clknet_1_1__leaf_net368));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net931 (.A(net931),
    .X(clknet_0_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_0__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net931 (.A(clknet_0_net931),
    .X(clknet_1_1__leaf_net931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net140 (.A(net140),
    .X(clknet_0_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_0__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net140 (.A(clknet_0_net140),
    .X(clknet_1_1__leaf_net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net153 (.A(net153),
    .X(clknet_0_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_0__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net153 (.A(clknet_0_net153),
    .X(clknet_1_1__leaf_net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net144 (.A(net144),
    .X(clknet_0_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_0__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net144 (.A(clknet_0_net144),
    .X(clknet_1_1__leaf_net144));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net145 (.A(net145),
    .X(clknet_0_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_0__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net145 (.A(clknet_0_net145),
    .X(clknet_1_1__leaf_net145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net142 (.A(net142),
    .X(clknet_0_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_0__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net142 (.A(clknet_0_net142),
    .X(clknet_1_1__leaf_net142));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net141 (.A(net141),
    .X(clknet_0_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_0__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net141 (.A(clknet_0_net141),
    .X(clknet_1_1__leaf_net141));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net128 (.A(net128),
    .X(clknet_0_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_0__leaf_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net128 (.A(clknet_0_net128),
    .X(clknet_1_1__leaf_net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net121 (.A(net121),
    .X(clknet_0_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net121 (.A(clknet_0_net121),
    .X(clknet_1_0__leaf_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net121 (.A(clknet_0_net121),
    .X(clknet_1_1__leaf_net121));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net998 (.A(net998),
    .X(clknet_0_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net998 (.A(clknet_0_net998),
    .X(clknet_1_0__leaf_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net998 (.A(clknet_0_net998),
    .X(clknet_1_1__leaf_net998));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net895 (.A(net895),
    .X(clknet_0_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_0__leaf_net895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net895 (.A(clknet_0_net895),
    .X(clknet_1_1__leaf_net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net882),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net591),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net252),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net826),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net426),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net431),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net231),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net111),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net747),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net893),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net740),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net239),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net939),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net600),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net916),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net869),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net905),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net178),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net305),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net870),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net41),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net584),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net595),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net868),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net642),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net783),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net392),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net738),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net874),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net842),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net876),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net523),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net245),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net813),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net176),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net809),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net787),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net589),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net681),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net709),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net599),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net872),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net438),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net805),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net394),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net969),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net39),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net40),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net755),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net391),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net795),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net31),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net921),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net458),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net810),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net597),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net912),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net867),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net925),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net875),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net918),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net643),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net853),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net244),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net314),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net777),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net403),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net786),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net591),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net234),
    .X(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_SCD (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_c154_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge804_C_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c290_B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c177_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c174_C (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_c155_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_S1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_D_N (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_SCE (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c163_C (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_c156_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c178_B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c162_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_c159_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_DE (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_S1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c335_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c334_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c226_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c201_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_c200_X (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c617_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_c240_Q (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_D (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge778_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge761_D (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c401_SET_B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c298_C1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A3 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_C1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_c270_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_S1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c277_B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_c276_X (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge861_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_S0 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c285_A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c284_A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c283_D_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_C (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_c278_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_SCE (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c442_B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c346_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c326_C (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_DE (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c452_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_Q (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_SCD (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c66_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_Q_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_S1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c633_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_SET_B (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_c359_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_S0 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c378_B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c375_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_c374_X (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_RESET_B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_D (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_DE (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_c417_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge780_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c65_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c45_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_c44_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_A0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_c438_X (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_D (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_SCE (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_SCD (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCE (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_SCD (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_C (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_c445_X (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_SCE (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_SCD (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c460_S0 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_RESET_B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c455_B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_c453_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_A0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_S0 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_A3 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_c463_X (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge840_A3 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_SCE (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_S0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_c465_X (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_SCE (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_A1 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge847_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge838_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c474_B (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c470_C (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_c469_X (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_SET_B (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_SCE (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_SCE (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c478_A3 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_c475_X (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_SCD (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c599_B (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_SCE (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c501_S0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c495_C (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_c482_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge848_A3 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_SCD (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_X (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_SET_B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_D_N (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c82_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_c75_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_A0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_Q_N (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_SCE (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_SCD (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_SCD (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c561_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_c554_X (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_Q (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_A2 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_C (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_c568_X (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_D (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c725_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_A3 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_SCD (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_A3 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_A3 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c726_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c626_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c613_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c612_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c607_S1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_Q (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_SCE (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge764_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c746_S0 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c632_B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_X (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_SCE (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_c95_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_X (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_c557_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_Q (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge762_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_Q (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c83_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_c473_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_net897_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_GCLK (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_c593_X (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_RESET_B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c130_C1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_SET_B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c121_B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c115_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c114_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_c113_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_Q (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_S0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_c287_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge904_Q (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c242_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_c196_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_Q_N (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_c189_S1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_Q (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c87_D1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c510_B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c484_C (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_A3 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_c32_B (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_SCE (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_SCE (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_SCE (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_SET_B (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_c489_X (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_X (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c255_D1 (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c120_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c112_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c110_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c96_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c104_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c103_C_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_B (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_c364_D_N (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c171_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge765_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge867_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge876_GATE_N (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge907_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge911_GATE (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge914_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge916_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_X (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c433_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c538_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c555_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge812_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge869_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_GATE (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge897_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s942_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c324_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_CLK_N (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge767_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge779_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_X (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s936_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c570_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c671_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c672_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge757_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge872_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge913_GATE (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s937_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c458_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c583_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c598_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge770_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge796_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge802_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge807_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_GATE (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s927_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s934_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c712_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c721_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c753_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge915_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s939_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c606_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c610_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c634_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c637_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge790_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge871_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge889_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge899_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s922_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s931_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s943_GATE_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c213_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c365_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c370_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c372_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge791_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge853_CLK_N (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge917_CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_X (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c125_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c127_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c131_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c219_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_CLK_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge888_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge902_CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge906_GATE (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge909_GATE_N (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_X (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c388_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge815_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge832_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge833_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge912_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s935_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s938_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S0 (.DIODE(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_S0 (.DIODE(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge852_S1 (.DIODE(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_S0 (.DIODE(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net503_X (.DIODE(clknet_1_0__leaf_net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_c511_A (.DIODE(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_c519_S1 (.DIODE(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_A3 (.DIODE(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge859_S1 (.DIODE(clknet_1_0__leaf_net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net365_X (.DIODE(clknet_1_0__leaf_net365));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
