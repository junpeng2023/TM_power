module netlist_0 (clk,
    in0,
    in1,
    in10,
    in11,
    in12,
    in13,
    in14,
    in15,
    in16,
    in17,
    in18,
    in19,
    in2,
    in20,
    in21,
    in22,
    in23,
    in24,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out0,
    out1,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
    out16,
    out17,
    out18,
    out19,
    out2,
    out20,
    out21,
    out22,
    out23,
    out24,
    out3,
    out4,
    out5,
    out6,
    out7,
    out8,
    out9,
    rst);
 input clk;
 input in0;
 input in1;
 input in10;
 input in11;
 input in12;
 input in13;
 input in14;
 input in15;
 input in16;
 input in17;
 input in18;
 input in19;
 input in2;
 input in20;
 input in21;
 input in22;
 input in23;
 input in24;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out0;
 output out1;
 output out10;
 output out11;
 output out12;
 output out13;
 output out14;
 output out15;
 output out16;
 output out17;
 output out18;
 output out19;
 output out2;
 output out20;
 output out21;
 output out22;
 output out23;
 output out24;
 output out3;
 output out4;
 output out5;
 output out6;
 output out7;
 output out8;
 output out9;
 input rst;

 wire net0;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net648;
 wire net754;
 wire net815;
 wire net911;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_0_net945;
 wire clknet_1_0__leaf_net945;
 wire clknet_1_1__leaf_net945;
 wire clknet_0_net260;
 wire clknet_1_0__leaf_net260;
 wire clknet_1_1__leaf_net260;
 wire clknet_0_net255;
 wire clknet_1_0__leaf_net255;
 wire clknet_1_1__leaf_net255;
 wire clknet_0_net944;
 wire clknet_1_0__leaf_net944;
 wire clknet_1_1__leaf_net944;
 wire clknet_0_net794;
 wire clknet_1_0__leaf_net794;
 wire clknet_1_1__leaf_net794;
 wire clknet_0_net745;
 wire clknet_1_0__leaf_net745;
 wire clknet_1_1__leaf_net745;
 wire clknet_0_net302;
 wire clknet_1_0__leaf_net302;
 wire clknet_1_1__leaf_net302;
 wire clknet_0_net301;
 wire clknet_1_0__leaf_net301;
 wire clknet_1_1__leaf_net301;
 wire clknet_0_net321;
 wire clknet_1_0__leaf_net321;
 wire clknet_1_1__leaf_net321;
 wire clknet_0_net307;
 wire clknet_1_0__leaf_net307;
 wire clknet_1_1__leaf_net307;
 wire clknet_0_net310;
 wire clknet_1_0__leaf_net310;
 wire clknet_1_1__leaf_net310;
 wire clknet_0_net759;
 wire clknet_1_0__leaf_net759;
 wire clknet_1_1__leaf_net759;
 wire clknet_0_net138;
 wire clknet_1_0__leaf_net138;
 wire clknet_1_1__leaf_net138;
 wire clknet_0_net135;
 wire clknet_1_0__leaf_net135;
 wire clknet_1_1__leaf_net135;
 wire clknet_0_net157;
 wire clknet_1_0__leaf_net157;
 wire clknet_1_1__leaf_net157;
 wire clknet_0_net178;
 wire clknet_1_0__leaf_net178;
 wire clknet_1_1__leaf_net178;
 wire clknet_0_net196;
 wire clknet_1_0__leaf_net196;
 wire clknet_1_1__leaf_net196;
 wire clknet_0_net164;
 wire clknet_1_0__leaf_net164;
 wire clknet_1_1__leaf_net164;
 wire clknet_0_net943;
 wire clknet_1_0__leaf_net943;
 wire clknet_1_1__leaf_net943;
 wire clknet_0_net33;
 wire clknet_1_0__leaf_net33;
 wire clknet_1_1__leaf_net33;
 wire clknet_0_net924;
 wire clknet_1_0__leaf_net924;
 wire clknet_1_1__leaf_net924;
 wire clknet_0_net585;
 wire clknet_1_0__leaf_net585;
 wire clknet_1_1__leaf_net585;
 wire clknet_0_net923;
 wire clknet_1_0__leaf_net923;
 wire clknet_1_1__leaf_net923;
 wire clknet_0_net655;
 wire clknet_1_0__leaf_net655;
 wire clknet_1_1__leaf_net655;
 wire clknet_0_net666;
 wire clknet_1_0__leaf_net666;
 wire clknet_1_1__leaf_net666;
 wire clknet_0_net660;
 wire clknet_1_0__leaf_net660;
 wire clknet_1_1__leaf_net660;
 wire clknet_0_net657;
 wire clknet_1_0__leaf_net657;
 wire clknet_1_1__leaf_net657;
 wire clknet_0_net652;
 wire clknet_1_0__leaf_net652;
 wire clknet_1_1__leaf_net652;
 wire clknet_0_net574;
 wire clknet_1_0__leaf_net574;
 wire clknet_1_1__leaf_net574;
 wire clknet_0_net898;
 wire clknet_1_0__leaf_net898;
 wire clknet_1_1__leaf_net898;
 wire clknet_0_net686;
 wire clknet_1_0__leaf_net686;
 wire clknet_1_1__leaf_net686;
 wire clknet_0_net922;
 wire clknet_1_0__leaf_net922;
 wire clknet_1_1__leaf_net922;
 wire clknet_0_net514;
 wire clknet_1_0__leaf_net514;
 wire clknet_1_1__leaf_net514;
 wire clknet_0_net523;
 wire clknet_1_0__leaf_net523;
 wire clknet_1_1__leaf_net523;
 wire clknet_0_net532;
 wire clknet_1_0__leaf_net532;
 wire clknet_1_1__leaf_net532;
 wire clknet_0_net528;
 wire clknet_1_0__leaf_net528;
 wire clknet_1_1__leaf_net528;
 wire clknet_0_net525;
 wire clknet_1_0__leaf_net525;
 wire clknet_1_1__leaf_net525;
 wire clknet_0_net516;
 wire clknet_1_0__leaf_net516;
 wire clknet_1_1__leaf_net516;
 wire clknet_0_net515;
 wire clknet_1_0__leaf_net515;
 wire clknet_1_1__leaf_net515;
 wire clknet_0_net413;
 wire clknet_1_0__leaf_net413;
 wire clknet_1_1__leaf_net413;
 wire clknet_0_net421;
 wire clknet_1_0__leaf_net421;
 wire clknet_1_1__leaf_net421;
 wire clknet_0_net414;
 wire clknet_1_0__leaf_net414;
 wire clknet_1_1__leaf_net414;
 wire clknet_0_net419;
 wire clknet_1_0__leaf_net419;
 wire clknet_1_1__leaf_net419;
 wire clknet_0_net415;
 wire clknet_1_0__leaf_net415;
 wire clknet_1_1__leaf_net415;
 wire clknet_0_net901;
 wire clknet_1_0__leaf_net901;
 wire clknet_1_1__leaf_net901;
 wire clknet_0_net439;
 wire clknet_1_0__leaf_net439;
 wire clknet_1_1__leaf_net439;
 wire clknet_0_net448;
 wire clknet_1_0__leaf_net448;
 wire clknet_1_1__leaf_net448;
 wire clknet_0_net445;
 wire clknet_1_0__leaf_net445;
 wire clknet_1_1__leaf_net445;
 wire clknet_0_net440;
 wire clknet_1_0__leaf_net440;
 wire clknet_1_1__leaf_net440;
 wire clknet_0_net441;
 wire clknet_1_0__leaf_net441;
 wire clknet_1_1__leaf_net441;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;

 sky130_fd_sc_hd__and2_1 c100 (.A(net79),
    .B(net77),
    .X(net80));
 sky130_fd_sc_hd__and2_1 c101 (.A(net78),
    .B(net77),
    .X(net81));
 sky130_fd_sc_hd__and3_1 c102 (.A(net72),
    .B(net80),
    .C(net81),
    .X(net82));
 sky130_fd_sc_hd__and2_0 c103 (.A(net81),
    .B(net77),
    .X(net83));
 sky130_fd_sc_hd__a2111o_1 c104 (.A1(net83),
    .A2(net82),
    .B1(net81),
    .C1(net80),
    .D1(net72),
    .X(net84));
 sky130_fd_sc_hd__and2_1 c105 (.A(net80),
    .B(net906),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 c106 (.A0(net85),
    .A1(net72),
    .A2(net80),
    .A3(net74),
    .S0(net78),
    .S1(net81),
    .X(net86));
 sky130_fd_sc_hd__buf_1 c107 (.A(net779),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 c108 (.A0(net78),
    .A1(net85),
    .A2(net87),
    .A3(net72),
    .S0(net81),
    .S1(net906),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 c109 (.A0(net88),
    .A1(net87),
    .A2(net85),
    .A3(net78),
    .S0(net79),
    .S1(net77),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 c110 (.A(net87),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 c111 (.A(net90),
    .X(net91));
 sky130_fd_sc_hd__buf_1 c112 (.X(net92));
 sky130_fd_sc_hd__and2_0 c113 (.A(net92),
    .B(net90),
    .X(net93));
 sky130_fd_sc_hd__and2_0 c114 (.A(net92),
    .B(net87),
    .X(net94));
 sky130_fd_sc_hd__and2_0 c115 (.A(net93),
    .B(net90),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 c116 (.A(net757),
    .X(net96));
 sky130_fd_sc_hd__and2_1 c117 (.A(net96),
    .B(net90),
    .X(net97));
 sky130_fd_sc_hd__and2_1 c118 (.A(net94),
    .B(net93),
    .X(net98));
 sky130_fd_sc_hd__buf_1 c119 (.A(net825),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 c120 (.A(net812),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 c121 (.A(net827),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 c122 (.A(net825),
    .X(net102));
 sky130_fd_sc_hd__and3_1 c123 (.A(net102),
    .B(net99),
    .C(net98),
    .X(net103));
 sky130_fd_sc_hd__and2_0 c124 (.A(net91),
    .B(net97),
    .X(net104));
 sky130_fd_sc_hd__and2_0 c125 (.A(net90),
    .B(net99),
    .X(net105));
 sky130_fd_sc_hd__and2_1 c126 (.A(net99),
    .B(net893),
    .X(net106));
 sky130_fd_sc_hd__and3_1 c127 (.A(net104),
    .B(net106),
    .C(net97),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 c128 (.A0(net106),
    .A1(net98),
    .A2(net102),
    .A3(net99),
    .S0(net97),
    .S1(net1067),
    .X(net108));
 sky130_fd_sc_hd__and3_1 c129 (.A(net97),
    .B(net106),
    .C(net893),
    .X(net109));
 sky130_fd_sc_hd__and3_1 c130 (.A(net105),
    .B(net106),
    .C(net918),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 c131 (.A0(net110),
    .A1(net100),
    .A2(net106),
    .A3(net98),
    .S0(net90),
    .S1(net1076),
    .X(net111));
 sky130_fd_sc_hd__and2_2 c132 (.A(net978),
    .B(net961),
    .X(net112));
 sky130_fd_sc_hd__and2_2 c133 (.A(net112),
    .B(net979),
    .X(net113));
 sky130_fd_sc_hd__and2_0 c134 (.A(net113),
    .B(net112),
    .X(net114));
 sky130_fd_sc_hd__and2_0 c135 (.A(net112),
    .B(net959),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 c136 (.A(net880),
    .X(net116));
 sky130_fd_sc_hd__and2_1 c137 (.A(net116),
    .B(net112),
    .X(net117));
 sky130_fd_sc_hd__and2_1 c138 (.A(net112),
    .B(net974),
    .X(net118));
 sky130_fd_sc_hd__and2_0 c139 (.A(net115),
    .B(net975),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 c140 (.A(net880),
    .X(net120));
 sky130_fd_sc_hd__and3_1 c141 (.A(net120),
    .B(net977),
    .C(net112),
    .X(net121));
 sky130_fd_sc_hd__and2_2 c142 (.A(net973),
    .B(net116),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 c143 (.A(net880),
    .X(net123));
 sky130_fd_sc_hd__and3_1 c144 (.A(net118),
    .B(net120),
    .C(net113),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 c145 (.A(net880),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 c146 (.A0(net125),
    .A1(net115),
    .A2(net123),
    .A3(net122),
    .S0(net113),
    .S1(net112),
    .X(net126));
 sky130_fd_sc_hd__and2_2 c147 (.A(net123),
    .B(net113),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 c148 (.A(net822),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 c149 (.A(net936),
    .X(net129));
 sky130_fd_sc_hd__and3_1 c150 (.A(net113),
    .B(net125),
    .C(net129),
    .X(net130));
 sky130_fd_sc_hd__buf_12 c151 (.A(net933),
    .X(net131));
 sky130_fd_sc_hd__and3_1 c152 (.A(net117),
    .B(net131),
    .C(net128),
    .X(net132));
 sky130_fd_sc_hd__buf_1 c153 (.A(net938),
    .X(net133));
 sky130_fd_sc_hd__buf_1 c154 (.A(net129),
    .X(net134));
 sky130_fd_sc_hd__buf_1 c155 (.A(clknet_1_0__leaf_net759),
    .X(net135));
 sky130_fd_sc_hd__and2_0 c156 (.A(net134),
    .B(net133),
    .X(net136));
 sky130_fd_sc_hd__buf_1 c157 (.A(net134),
    .X(net137));
 sky130_fd_sc_hd__buf_1 c158 (.A(clknet_1_1__leaf_net759),
    .X(net138));
 sky130_fd_sc_hd__and2_1 c159 (.A(net137),
    .B(net133),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 c160 (.A(net773),
    .X(net140));
 sky130_fd_sc_hd__and2_0 c161 (.A(clknet_1_1__leaf_net138),
    .B(net754),
    .X(net141));
 sky130_fd_sc_hd__and2_1 c162 (.A(net134),
    .B(net137),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 c163 (.X(net143));
 sky130_fd_sc_hd__and2_4 c164 (.A(net134),
    .B(net137),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 c165 (.A(net774),
    .X(net145));
 sky130_fd_sc_hd__and2_1 c166 (.A(net972),
    .B(net137),
    .X(net146));
 sky130_fd_sc_hd__buf_1 c167 (.A(net786),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 c168 (.A(net954),
    .X(net148));
 sky130_fd_sc_hd__buf_1 c169 (.A(net792),
    .X(net149));
 sky130_fd_sc_hd__and3_1 c170 (.A(net147),
    .B(net149),
    .C(net965),
    .X(net150));
 sky130_fd_sc_hd__and3_1 c171 (.A(net149),
    .B(net147),
    .C(net150),
    .X(net151));
 sky130_fd_sc_hd__a2111o_1 c172 (.A1(net140),
    .A2(net147),
    .B1(net149),
    .C1(net150),
    .D1(net144),
    .X(net152));
 sky130_fd_sc_hd__and3_1 c173 (.A(net148),
    .B(net150),
    .C(net871),
    .X(net153));
 sky130_fd_sc_hd__and3_1 c174 (.A(net150),
    .B(net153),
    .C(net1026),
    .X(net154));
 sky130_fd_sc_hd__or4bb_1 c175 (.A(net136),
    .B(net1027),
    .C_N(net150),
    .D_N(net144),
    .X(net155));
 sky130_fd_sc_hd__and2_0 c176 (.A(net967),
    .B(net36),
    .X(net156));
 sky130_fd_sc_hd__buf_1 c177 (.A(clknet_1_1__leaf_net135),
    .X(net157));
 sky130_fd_sc_hd__and2_1 c178 (.A(net133),
    .B(net871),
    .X(net158));
 sky130_fd_sc_hd__buf_1 c179 (.A(net761),
    .X(net159));
 sky130_fd_sc_hd__and2_0 c180 (.A(clknet_1_0__leaf_net157),
    .B(net158),
    .X(net160));
 sky130_fd_sc_hd__and2_0 c181 (.A(net24),
    .B(net158),
    .X(net161));
 sky130_fd_sc_hd__and2_0 c182 (.A(net151),
    .B(net158),
    .X(net162));
 sky130_fd_sc_hd__and2_1 c183 (.A(net159),
    .B(net24),
    .X(net163));
 sky130_fd_sc_hd__and2_0 c184 (.A(net160),
    .B(net163),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 c185 (.A(net761),
    .X(net165));
 sky130_fd_sc_hd__and2_1 c186 (.A(net165),
    .B(net159),
    .X(net166));
 sky130_fd_sc_hd__and3_1 c187 (.A(net161),
    .B(net166),
    .C(clknet_1_0__leaf_net164),
    .X(net167));
 sky130_fd_sc_hd__and2_0 c188 (.A(net158),
    .B(net166),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 c189 (.A(net856),
    .X(net169));
 sky130_fd_sc_hd__and2_0 c190 (.A(net169),
    .B(net873),
    .X(net170));
 sky130_fd_sc_hd__and2_0 c191 (.A(net156),
    .B(net159),
    .X(net171));
 sky130_fd_sc_hd__buf_1 c192 (.A(net855),
    .X(net172));
 sky130_fd_sc_hd__and3_1 c193 (.A(net168),
    .B(net171),
    .C(net172),
    .X(net173));
 sky130_fd_sc_hd__and3_1 c194 (.A(net172),
    .B(net163),
    .C(net168),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 c195 (.A(net1044),
    .X(net175));
 sky130_fd_sc_hd__and3_1 c196 (.A(net175),
    .B(net174),
    .C(net168),
    .X(net176));
 sky130_fd_sc_hd__and3_1 c197 (.A(net170),
    .B(net166),
    .C(net872),
    .X(net177));
 sky130_fd_sc_hd__buf_1 c198 (.A(clknet_1_1__leaf_net157),
    .X(net178));
 sky130_fd_sc_hd__buf_1 c199 (.A(clknet_1_0__leaf_net178),
    .X(net179));
 sky130_fd_sc_hd__buf_1 c200 (.A(net891),
    .X(net180));
 sky130_fd_sc_hd__and2_1 c201 (.A(net180),
    .B(net891),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 c202 (.A(net760),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 c203 (.A(net760),
    .X(net183));
 sky130_fd_sc_hd__and2_1 c204 (.A(net183),
    .B(net177),
    .X(net184));
 sky130_fd_sc_hd__and2_0 c205 (.A(net181),
    .B(net183),
    .X(net185));
 sky130_fd_sc_hd__buf_1 c206 (.A(net818),
    .X(net186));
 sky130_fd_sc_hd__buf_1 c207 (.A(net782),
    .X(net187));
 sky130_fd_sc_hd__and2_0 c208 (.A(net186),
    .B(net181),
    .X(net188));
 sky130_fd_sc_hd__and3_1 c209 (.A(net183),
    .B(net186),
    .C(clknet_1_1__leaf_net178),
    .X(net189));
 sky130_fd_sc_hd__and2_0 c210 (.A(net186),
    .B(net182),
    .X(net190));
 sky130_fd_sc_hd__and2_1 c211 (.A(net187),
    .B(net181),
    .X(net191));
 sky130_fd_sc_hd__mux4_1 c212 (.A0(net188),
    .A1(clknet_1_0__leaf_net178),
    .A2(net191),
    .A3(net56),
    .S0(net57),
    .S1(net186),
    .X(net192));
 sky130_fd_sc_hd__and3_1 c213 (.A(net182),
    .B(net187),
    .C(net886),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 c214 (.A(net806),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 c215 (.A(net929),
    .X(net195));
 sky130_fd_sc_hd__or4bb_1 c216 (.A(clknet_1_1__leaf_net178),
    .B(net194),
    .C_N(net190),
    .D_N(net195),
    .X(net196));
 sky130_fd_sc_hd__and2_0 c217 (.A(net195),
    .B(net193),
    .X(net197));
 sky130_fd_sc_hd__sdfrbp_1 c218 (.CLK(clknet_4_11_0_clk),
    .D(net190),
    .RESET_B(clknet_1_1__leaf_net196),
    .SCD(net197),
    .SCE(net183),
    .Q(net199),
    .Q_N(net198));
 sky130_fd_sc_hd__or4bb_1 c219 (.A(net191),
    .B(net197),
    .C_N(net183),
    .D_N(clknet_1_0__leaf_net196),
    .X(net200));
 sky130_fd_sc_hd__and2_0 c220 (.A(net199),
    .B(net180),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 c221 (.A(net906),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 c222 (.A(net767),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 c223 (.A(net202),
    .X(net204));
 sky130_fd_sc_hd__and2_2 c224 (.A(net204),
    .B(net203),
    .X(net205));
 sky130_fd_sc_hd__and2_0 c225 (.A(net87),
    .B(net202),
    .X(net206));
 sky130_fd_sc_hd__and2_0 c226 (.A(net180),
    .B(net203),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 c227 (.A(net766),
    .X(net208));
 sky130_fd_sc_hd__and2_1 c228 (.A(net206),
    .B(net202),
    .X(net209));
 sky130_fd_sc_hd__dfbbn_1 c229 (.CLK_N(clknet_4_10_0_clk),
    .D(net209),
    .RESET_B(net206),
    .SET_B(net205),
    .Q(net211),
    .Q_N(net210));
 sky130_fd_sc_hd__buf_1 c230 (.A(net796),
    .X(net212));
 sky130_fd_sc_hd__dfbbp_1 c231 (.CLK(clknet_4_9_0_clk),
    .D(net212),
    .RESET_B(net205),
    .SET_B(net209),
    .Q(net214),
    .Q_N(net213));
 sky130_fd_sc_hd__clkbuf_1 c232 (.A(net823),
    .X(net215));
 sky130_fd_sc_hd__sdfxbp_1 c233 (.CLK(clknet_4_9_0_clk),
    .D(net215),
    .SCD(net205),
    .SCE(net213),
    .Q(net217),
    .Q_N(net216));
 sky130_fd_sc_hd__and2_0 c234 (.A(net203),
    .B(net201),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 c235 (.A(net949),
    .X(net219));
 sky130_fd_sc_hd__and2_0 c236 (.A(net202),
    .B(net219),
    .X(net220));
 sky130_fd_sc_hd__and3_1 c237 (.A(net214),
    .B(net205),
    .C(net209),
    .X(net221));
 sky130_fd_sc_hd__sdfxbp_1 c238 (.CLK(clknet_4_8_0_clk),
    .D(net218),
    .SCD(net202),
    .SCE(net1074),
    .Q(net223),
    .Q_N(net222));
 sky130_fd_sc_hd__and3_1 c239 (.A(net219),
    .B(net207),
    .C(net1081),
    .X(net224));
 sky130_fd_sc_hd__and3_1 c240 (.A(net220),
    .B(net1020),
    .C(net224),
    .X(net225));
 sky130_fd_sc_hd__sdfxtp_1 c241 (.CLK(clknet_4_9_0_clk),
    .D(net1032),
    .SCD(net224),
    .SCE(net1071),
    .Q(net226));
 sky130_fd_sc_hd__and2_0 c242 (.A(net92),
    .B(net885),
    .X(net227));
 sky130_fd_sc_hd__and2_0 c243 (.A(net227),
    .B(net92),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 c244 (.A(net749),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 c245 (.A(net211),
    .X(net230));
 sky130_fd_sc_hd__and2_2 c246 (.A(net229),
    .B(net228),
    .X(net231));
 sky130_fd_sc_hd__sdfxtp_1 c247 (.CLK(clknet_4_10_0_clk),
    .D(net1041),
    .SCD(net231),
    .SCE(net1043),
    .Q(net232));
 sky130_fd_sc_hd__sdfxtp_1 c248 (.CLK(clknet_4_10_0_clk),
    .D(net228),
    .SCD(net231),
    .SCE(net1035),
    .Q(net233));
 sky130_fd_sc_hd__clkbuf_1 c249 (.A(net749),
    .X(net234));
 sky130_fd_sc_hd__and2_1 c25 (.A(net970),
    .B(net815),
    .X(net0));
 sky130_fd_sc_hd__clkbuf_1 c250 (.A(net798),
    .X(net235));
 sky130_fd_sc_hd__and2_0 c251 (.A(net235),
    .B(net232),
    .X(net236));
 sky130_fd_sc_hd__dfbbn_1 c252 (.CLK_N(clknet_4_10_0_clk),
    .D(net232),
    .RESET_B(net229),
    .SET_B(net231),
    .Q(net238),
    .Q_N(net237));
 sky130_fd_sc_hd__buf_1 c253 (.A(net798),
    .X(net239));
 sky130_fd_sc_hd__and3_1 c254 (.A(net236),
    .B(net233),
    .C(net239),
    .X(net240));
 sky130_fd_sc_hd__and3_1 c255 (.A(net239),
    .B(net240),
    .C(net238),
    .X(net241));
 sky130_fd_sc_hd__and3_1 c256 (.A(net241),
    .B(net238),
    .C(net239),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 c257 (.A(net930),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 c258 (.A(net931),
    .X(net244));
 sky130_fd_sc_hd__or4bb_1 c259 (.A(net230),
    .B(net235),
    .C_N(net240),
    .D_N(net1035),
    .X(net245));
 sky130_fd_sc_hd__and3_1 c26 (.A(net0),
    .B(net648),
    .C(net976),
    .X(net1));
 sky130_fd_sc_hd__or4bb_1 c260 (.A(net234),
    .B(net245),
    .C_N(net1035),
    .D_N(net231),
    .X(net246));
 sky130_fd_sc_hd__and3_1 c261 (.A(net244),
    .B(net227),
    .C(net919),
    .X(net247));
 sky130_fd_sc_hd__and3_1 c262 (.A(net247),
    .B(net239),
    .C(net879),
    .X(net248));
 sky130_fd_sc_hd__mux4_1 c263 (.A0(net248),
    .A1(net234),
    .A2(net243),
    .A3(net241),
    .S0(net237),
    .S1(net231),
    .X(net249));
 sky130_fd_sc_hd__buf_12 c264 (.A(net131),
    .X(net250));
 sky130_fd_sc_hd__and2_0 c265 (.A(net133),
    .B(net250),
    .X(net251));
 sky130_fd_sc_hd__buf_2 c266 (.A(net734),
    .X(net252));
 sky130_fd_sc_hd__and2_4 c267 (.A(net252),
    .B(net250),
    .X(net253));
 sky130_fd_sc_hd__buf_1 c268 (.A(net733),
    .X(net254));
 sky130_fd_sc_hd__buf_1 c269 (.A(clknet_1_0__leaf_net945),
    .X(net255));
 sky130_fd_sc_hd__and2_0 c27 (.A(net971),
    .B(net960),
    .X(net2));
 sky130_fd_sc_hd__and2_0 c270 (.A(clknet_1_0__leaf_net255),
    .B(net254),
    .X(net256));
 sky130_fd_sc_hd__and3_4 c271 (.A(net250),
    .B(net254),
    .C(net252),
    .X(net257));
 sky130_fd_sc_hd__and3_1 c272 (.A(net251),
    .B(clknet_1_1__leaf_net255),
    .C(net250),
    .X(net258));
 sky130_fd_sc_hd__and2_0 c273 (.A(clknet_1_0__leaf_net255),
    .B(net257),
    .X(net259));
 sky130_fd_sc_hd__buf_1 c274 (.A(clknet_1_1__leaf_net945),
    .X(net260));
 sky130_fd_sc_hd__and3_1 c275 (.A(clknet_1_0__leaf_net260),
    .B(net257),
    .C(net254),
    .X(net261));
 sky130_fd_sc_hd__and3_1 c276 (.A(net261),
    .B(net257),
    .C(clknet_1_1__leaf_net260),
    .X(net262));
 sky130_fd_sc_hd__buf_1 c277 (.A(net953),
    .X(net263));
 sky130_fd_sc_hd__and3_4 c278 (.A(net257),
    .B(net253),
    .C(net263),
    .X(net264));
 sky130_fd_sc_hd__dfbbn_1 c279 (.CLK_N(clknet_4_0_0_clk),
    .D(net256),
    .RESET_B(net264),
    .SET_B(clknet_1_0__leaf_net260),
    .Q(net266),
    .Q_N(net265));
 sky130_fd_sc_hd__and3_1 c28 (.A(net8),
    .B(net971),
    .C(net0),
    .X(net3));
 sky130_fd_sc_hd__sdfrtn_1 c280 (.CLK_N(clknet_4_0_0_clk),
    .D(net254),
    .RESET_B(net1019),
    .SCD(net264),
    .SCE(net127),
    .Q(net267));
 sky130_fd_sc_hd__sdfbbn_1 c281 (.CLK_N(clknet_4_1_0_clk),
    .D(net1073),
    .RESET_B(net1029),
    .SCD(net1064),
    .SCE(net264),
    .SET_B(net996),
    .Q(net269),
    .Q_N(net268));
 sky130_fd_sc_hd__a2111o_1 c282 (.A1(net258),
    .A2(net269),
    .B1(net263),
    .C1(net994),
    .D1(net252),
    .X(net270));
 sky130_fd_sc_hd__dfbbp_1 c283 (.CLK(clknet_4_1_0_clk),
    .D(net269),
    .RESET_B(net264),
    .SET_B(net267),
    .Q(net271));
 sky130_fd_sc_hd__a2111o_1 c284 (.A1(net271),
    .A2(net268),
    .B1(net267),
    .C1(net995),
    .D1(net884),
    .X(net272));
 sky130_fd_sc_hd__sdfbbn_1 c285 (.CLK_N(clknet_4_1_0_clk),
    .D(net132),
    .RESET_B(net994),
    .SCD(net250),
    .SCE(net1077),
    .SET_B(net908),
    .Q(net273));
 sky130_fd_sc_hd__buf_1 c286 (.A(net771),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 c287 (.A(net274),
    .X(net275));
 sky130_fd_sc_hd__and2_1 c288 (.A(net274),
    .B(net252),
    .X(net276));
 sky130_fd_sc_hd__and3_1 c289 (.A(net276),
    .B(net275),
    .C(net19),
    .X(net277));
 sky130_fd_sc_hd__and2_0 c29 (.A(net970),
    .B(net971),
    .X(net4));
 sky130_fd_sc_hd__and2_0 c290 (.A(net277),
    .B(net276),
    .X(net278));
 sky130_fd_sc_hd__buf_1 c291 (.A(net771),
    .X(net279));
 sky130_fd_sc_hd__and2_0 c292 (.A(net277),
    .B(net279),
    .X(net280));
 sky130_fd_sc_hd__and2_1 c293 (.A(net276),
    .B(net279),
    .X(net281));
 sky130_fd_sc_hd__and3_1 c294 (.A(net275),
    .B(net276),
    .C(net279),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 c295 (.A(net1080),
    .X(net283));
 sky130_fd_sc_hd__and2_1 c296 (.A(net279),
    .B(net283),
    .X(net284));
 sky130_fd_sc_hd__and2_2 c297 (.A(net282),
    .B(net281),
    .X(net285));
 sky130_fd_sc_hd__buf_1 c298 (.A(net940),
    .X(net286));
 sky130_fd_sc_hd__and3_1 c299 (.A(net139),
    .B(net285),
    .C(net279),
    .X(net287));
 sky130_fd_sc_hd__or4bb_2 c30 (.A(net4),
    .B(net968),
    .C_N(net3),
    .D_N(net971),
    .X(net5));
 sky130_fd_sc_hd__sdfxbp_1 c300 (.CLK(clknet_4_1_0_clk),
    .D(net283),
    .SCD(net278),
    .SCE(net284),
    .Q(net289),
    .Q_N(net288));
 sky130_fd_sc_hd__sdfxbp_1 c301 (.CLK(clknet_4_3_0_clk),
    .D(net280),
    .SCD(net286),
    .SCE(net277),
    .Q(net291),
    .Q_N(net290));
 sky130_fd_sc_hd__or4bb_1 c302 (.A(net284),
    .B(net1060),
    .C_N(net279),
    .D_N(net286),
    .X(net292));
 sky130_fd_sc_hd__sdfbbp_1 c303 (.CLK(clknet_4_0_0_clk),
    .D(net292),
    .RESET_B(net280),
    .SCD(net276),
    .SCE(net285),
    .SET_B(net284),
    .Q(net294),
    .Q_N(net293));
 sky130_fd_sc_hd__and3_1 c304 (.A(net294),
    .B(net284),
    .C(net275),
    .X(net295));
 sky130_fd_sc_hd__a2111o_1 c305 (.A1(net274),
    .A2(net286),
    .B1(net288),
    .C1(net293),
    .D1(net276),
    .X(net296));
 sky130_fd_sc_hd__and3_1 c306 (.A(net278),
    .B(net294),
    .C(net295),
    .X(net297));
 sky130_fd_sc_hd__a2111o_1 c307 (.A1(net296),
    .A2(net290),
    .B1(net293),
    .C1(net145),
    .D1(net1069),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 c308 (.A(net177),
    .X(net299));
 sky130_fd_sc_hd__buf_1 c309 (.A(net295),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 c31 (.A(net756),
    .X(net6));
 sky130_fd_sc_hd__buf_1 c310 (.A(clknet_1_1__leaf_net745),
    .X(net301));
 sky130_fd_sc_hd__buf_1 c311 (.A(clknet_1_0__leaf_net745),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 c312 (.A(net889),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 c313 (.A(net781),
    .X(net304));
 sky130_fd_sc_hd__and2_1 c314 (.A(net303),
    .B(net892),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 c315 (.A(net832),
    .X(net306));
 sky130_fd_sc_hd__and2_0 c316 (.A(clknet_1_1__leaf_net301),
    .B(net305),
    .X(net307));
 sky130_fd_sc_hd__and2_0 c317 (.A(net306),
    .B(clknet_1_0__leaf_net307),
    .X(net308));
 sky130_fd_sc_hd__buf_1 c318 (.A(clknet_1_0__leaf_net794),
    .X(net309));
 sky130_fd_sc_hd__and2_0 c319 (.A(clknet_1_0__leaf_net307),
    .B(net305),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 c32 (.A(net1065),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 c320 (.A(net952),
    .X(net311));
 sky130_fd_sc_hd__and3_1 c321 (.A(net309),
    .B(net303),
    .C(clknet_1_0__leaf_net301),
    .X(net312));
 sky130_fd_sc_hd__buf_1 c322 (.A(net950),
    .X(net313));
 sky130_fd_sc_hd__and2_0 c323 (.A(net304),
    .B(net313),
    .X(net314));
 sky130_fd_sc_hd__and2_0 c324 (.A(clknet_1_1__leaf_net157),
    .B(clknet_1_1__leaf_net301),
    .X(net315));
 sky130_fd_sc_hd__sdfxtp_2 c325 (.CLK(clknet_4_3_0_clk),
    .D(net305),
    .SCD(net314),
    .SCE(clknet_1_0__leaf_net310),
    .Q(net316));
 sky130_fd_sc_hd__clkbuf_1 c326 (.A(net937),
    .X(net317));
 sky130_fd_sc_hd__or4bb_1 c327 (.A(net315),
    .B(net316),
    .C_N(net313),
    .D_N(net303),
    .X(net318));
 sky130_fd_sc_hd__or4bb_1 c328 (.A(net317),
    .B(net318),
    .C_N(net303),
    .D_N(net316),
    .X(net319));
 sky130_fd_sc_hd__or4bb_1 c329 (.A(net312),
    .B(net316),
    .C_N(net313),
    .D_N(net889),
    .X(net320));
 sky130_fd_sc_hd__and2_1 c33 (.A(net911),
    .B(net963),
    .X(net8));
 sky130_fd_sc_hd__buf_1 c330 (.A(net320),
    .X(net321));
 sky130_fd_sc_hd__buf_2 c331 (.X(net322));
 sky130_fd_sc_hd__and2_4 c332 (.A(net67),
    .B(net199),
    .X(net323));
 sky130_fd_sc_hd__and2_0 c333 (.A(net322),
    .B(net180),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 c334 (.A(net770),
    .X(net325));
 sky130_fd_sc_hd__buf_1 c335 (.A(net928),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 c336 (.A(net955),
    .X(net327));
 sky130_fd_sc_hd__and2_0 c337 (.A(net325),
    .B(net322),
    .X(net328));
 sky130_fd_sc_hd__and2_1 c338 (.A(net327),
    .B(net325),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 c339 (.A(net789),
    .X(net330));
 sky130_fd_sc_hd__and2_1 c34 (.A(net0),
    .B(net7),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 c340 (.A(net819),
    .X(net331));
 sky130_fd_sc_hd__and2_0 c341 (.A(net328),
    .B(net330),
    .X(net332));
 sky130_fd_sc_hd__and3_1 c342 (.A(net331),
    .B(net326),
    .C(net329),
    .X(net333));
 sky130_fd_sc_hd__and3_2 c343 (.A(net56),
    .B(net330),
    .C(net322),
    .X(net334));
 sky130_fd_sc_hd__and2_1 c344 (.A(net332),
    .B(net334),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 c345 (.A(net889),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 c346 (.A(net935),
    .X(net337));
 sky130_fd_sc_hd__and3_1 c347 (.A(net303),
    .B(net336),
    .C(net337),
    .X(net338));
 sky130_fd_sc_hd__and3_1 c348 (.A(net337),
    .B(net335),
    .C(net334),
    .X(net339));
 sky130_fd_sc_hd__mux4_1 c349 (.A0(net338),
    .A1(net333),
    .A2(net337),
    .A3(net335),
    .S0(net322),
    .S1(net323),
    .X(net340));
 sky130_fd_sc_hd__and3_1 c35 (.A(net3),
    .B(net9),
    .C(net8),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 c350 (.A(net942),
    .X(net341));
 sky130_fd_sc_hd__buf_6 c351 (.A(net993),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 c352 (.A(net226),
    .X(net343));
 sky130_fd_sc_hd__buf_1 c353 (.A(net343),
    .X(net344));
 sky130_fd_sc_hd__and2_4 c354 (.A(net342),
    .B(net226),
    .X(net345));
 sky130_fd_sc_hd__buf_6 c355 (.A(net345),
    .X(net346));
 sky130_fd_sc_hd__and2_0 c356 (.A(net344),
    .B(net345),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 c357 (.A(net755),
    .X(net348));
 sky130_fd_sc_hd__and2_0 c358 (.A(net344),
    .B(net334),
    .X(net349));
 sky130_fd_sc_hd__and2_0 c359 (.A(net345),
    .B(net346),
    .X(net350));
 sky130_fd_sc_hd__dfbbn_1 c36 (.CLK_N(clknet_4_0_0_clk),
    .D(net969),
    .RESET_B(net10),
    .SET_B(net9),
    .Q(net12),
    .Q_N(net11));
 sky130_fd_sc_hd__and2_0 c360 (.A(net348),
    .B(net322),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 c361 (.A(net755),
    .X(net352));
 sky130_fd_sc_hd__and2_1 c362 (.A(net343),
    .B(net352),
    .X(net353));
 sky130_fd_sc_hd__and2_1 c363 (.A(net351),
    .B(net344),
    .X(net354));
 sky130_fd_sc_hd__and2_0 c364 (.A(net311),
    .B(net344),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 c365 (.A(net797),
    .X(net356));
 sky130_fd_sc_hd__and2_4 c366 (.A(net346),
    .B(net348),
    .X(net357));
 sky130_fd_sc_hd__sdfxtp_1 c367 (.CLK(clknet_4_14_0_clk),
    .D(net356),
    .SCD(net357),
    .SCE(net354),
    .Q(net358));
 sky130_fd_sc_hd__clkbuf_1 c368 (.A(net1021),
    .X(net359));
 sky130_fd_sc_hd__or4bb_1 c369 (.A(net353),
    .B(net354),
    .C_N(net345),
    .D_N(net359),
    .X(net360));
 sky130_fd_sc_hd__and3_1 c37 (.A(net9),
    .B(net3),
    .C(net11),
    .X(net13));
 sky130_fd_sc_hd__and3_1 c370 (.A(net359),
    .B(net354),
    .C(net345),
    .X(net361));
 sky130_fd_sc_hd__sdfxtp_1 c371 (.CLK(clknet_4_12_0_clk),
    .D(net357),
    .SCD(net354),
    .SCE(net1050),
    .Q(net362));
 sky130_fd_sc_hd__and2_1 c372 (.A(net362),
    .B(net864),
    .X(net363));
 sky130_fd_sc_hd__sdfbbn_1 c373 (.CLK_N(clknet_4_12_0_clk),
    .D(net352),
    .RESET_B(net359),
    .SCD(net363),
    .SCE(net357),
    .SET_B(net344),
    .Q(net364));
 sky130_fd_sc_hd__clkbuf_2 c374 (.A(net920),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 c375 (.A(net365),
    .X(net366));
 sky130_fd_sc_hd__and2_1 c376 (.A(net365),
    .B(net920),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 c377 (.X(net368));
 sky130_fd_sc_hd__and2_1 c378 (.A(net366),
    .B(net368),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 c379 (.A(net753),
    .X(net370));
 sky130_fd_sc_hd__a2111o_1 c38 (.A1(net971),
    .A2(net12),
    .B1(net970),
    .C1(net5),
    .D1(net8),
    .X(net14));
 sky130_fd_sc_hd__dfbbn_1 c380 (.CLK_N(clknet_4_14_0_clk),
    .D(net1033),
    .RESET_B(net369),
    .SET_B(net365),
    .Q(net372),
    .Q_N(net371));
 sky130_fd_sc_hd__and2_2 c381 (.A(net372),
    .B(net365),
    .X(net373));
 sky130_fd_sc_hd__or4bb_1 c382 (.A(net334),
    .B(net369),
    .C_N(net371),
    .D_N(net373),
    .X(net374));
 sky130_fd_sc_hd__and2_1 c383 (.A(net370),
    .B(net1046),
    .X(net375));
 sky130_fd_sc_hd__and3_1 c384 (.A(net369),
    .B(net370),
    .C(net365),
    .X(net376));
 sky130_fd_sc_hd__dfbbn_1 c385 (.CLK_N(clknet_4_14_0_clk),
    .D(net375),
    .RESET_B(net357),
    .SET_B(net373),
    .Q(net378),
    .Q_N(net377));
 sky130_fd_sc_hd__and2_1 c386 (.A(net373),
    .B(net378),
    .X(net379));
 sky130_fd_sc_hd__sdfrtp_1 c387 (.CLK(clknet_4_14_0_clk),
    .D(net378),
    .RESET_B(net1047),
    .SCD(net373),
    .SCE(net1068),
    .Q(net380));
 sky130_fd_sc_hd__clkbuf_1 c388 (.A(net955),
    .X(net381));
 sky130_fd_sc_hd__and3_1 c389 (.A(net381),
    .B(net366),
    .C(net365),
    .X(net382));
 sky130_fd_sc_hd__and3_1 c39 (.A(net962),
    .B(net971),
    .C(net897),
    .X(net15));
 sky130_fd_sc_hd__sdfrtp_1 c390 (.CLK(clknet_4_14_0_clk),
    .D(net365),
    .RESET_B(net1055),
    .SCD(net372),
    .SCE(net375),
    .Q(net383));
 sky130_fd_sc_hd__clkbuf_1 c391 (.A(net948),
    .X(net384));
 sky130_fd_sc_hd__buf_1 c392 (.A(clknet_1_1__leaf_net943),
    .X(net385));
 sky130_fd_sc_hd__and3_1 c393 (.A(net385),
    .B(net380),
    .C(net377),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 c394 (.A(net935),
    .X(net387));
 sky130_fd_sc_hd__sdfrtp_1 c395 (.CLK(clknet_4_11_0_clk),
    .D(net386),
    .RESET_B(net1018),
    .SCD(net387),
    .SCE(net379),
    .Q(net388));
 sky130_fd_sc_hd__and2_2 c396 (.A(net273),
    .B(net252),
    .X(net389));
 sky130_fd_sc_hd__buf_1 c397 (.A(net389),
    .X(net390));
 sky130_fd_sc_hd__and2_1 c398 (.A(net252),
    .B(net389),
    .X(net391));
 sky130_fd_sc_hd__and2_1 c399 (.A(net389),
    .B(net390),
    .X(net392));
 sky130_fd_sc_hd__or4bb_1 c40 (.A(net1),
    .B(net13),
    .C_N(net3),
    .D_N(net9),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 c400 (.A(net739),
    .X(net393));
 sky130_fd_sc_hd__and3_1 c401 (.A(net393),
    .B(net390),
    .C(net391),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 c402 (.A(net932),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 c403 (.A(net958),
    .X(net396));
 sky130_fd_sc_hd__and2_1 c404 (.A(net396),
    .B(net390),
    .X(net397));
 sky130_fd_sc_hd__buf_1 c405 (.A(net1059),
    .X(net398));
 sky130_fd_sc_hd__and2_1 c406 (.A(net390),
    .B(net396),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 c407 (.A(net740),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 c408 (.A(net957),
    .X(net401));
 sky130_fd_sc_hd__and3_1 c409 (.A(net122),
    .B(net399),
    .C(net398),
    .X(net402));
 sky130_fd_sc_hd__or4bb_1 c41 (.A(net6),
    .B(net12),
    .C_N(net966),
    .D_N(net9),
    .X(net17));
 sky130_fd_sc_hd__a2111o_1 c410 (.A1(net392),
    .A2(net400),
    .B1(net398),
    .C1(net393),
    .D1(net252),
    .X(net403));
 sky130_fd_sc_hd__and3_1 c411 (.A(net398),
    .B(net390),
    .C(net878),
    .X(net404));
 sky130_fd_sc_hd__and3_1 c412 (.A(net398),
    .B(net393),
    .C(net878),
    .X(net405));
 sky130_fd_sc_hd__dfbbp_1 c413 (.CLK(clknet_4_4_0_clk),
    .D(net405),
    .RESET_B(net397),
    .SET_B(net393),
    .Q(net407),
    .Q_N(net406));
 sky130_fd_sc_hd__mux4_1 c414 (.A0(net395),
    .A1(net393),
    .A2(net406),
    .A3(net391),
    .S0(net389),
    .S1(net392),
    .X(net408));
 sky130_fd_sc_hd__sdfxbp_1 c415 (.CLK(clknet_4_4_0_clk),
    .D(net1078),
    .SCD(net404),
    .SCE(net1056),
    .Q(net410),
    .Q_N(net409));
 sky130_fd_sc_hd__and3_1 c416 (.A(net401),
    .B(net398),
    .C(net410),
    .X(net411));
 sky130_fd_sc_hd__mux4_1 c417 (.A0(net391),
    .A1(net411),
    .A2(net409),
    .A3(net398),
    .S0(net404),
    .S1(net1056),
    .X(net412));
 sky130_fd_sc_hd__buf_1 c418 (.A(clknet_1_0__leaf_net922),
    .X(net413));
 sky130_fd_sc_hd__buf_1 c419 (.A(clknet_1_0__leaf_net413),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 c42 (.A0(net17),
    .A1(net15),
    .A2(net12),
    .A3(net970),
    .S0(net5),
    .S1(net907),
    .X(net18));
 sky130_fd_sc_hd__buf_1 c420 (.A(clknet_1_0__leaf_net414),
    .X(net415));
 sky130_fd_sc_hd__buf_1 c421 (.A(net738),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 c422 (.A(net737),
    .X(net417));
 sky130_fd_sc_hd__and2_0 c423 (.A(net417),
    .B(clknet_1_0__leaf_net414),
    .X(net418));
 sky130_fd_sc_hd__buf_1 c424 (.A(clknet_1_1__leaf_net414),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 c425 (.A(net805),
    .X(net420));
 sky130_fd_sc_hd__and2_0 c426 (.A(clknet_1_1__leaf_net414),
    .B(clknet_1_0__leaf_net413),
    .X(net421));
 sky130_fd_sc_hd__buf_1 c427 (.A(net804),
    .X(net422));
 sky130_fd_sc_hd__buf_1 c428 (.A(net790),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 c429 (.A(net800),
    .X(net424));
 sky130_fd_sc_hd__sdfbbn_1 c43 (.CLK_N(clknet_4_2_0_clk),
    .D(net970),
    .RESET_B(net1054),
    .SCD(net5),
    .SCE(net897),
    .SET_B(net907),
    .Q(net20),
    .Q_N(net19));
 sky130_fd_sc_hd__or4bb_1 c430 (.A(net422),
    .B(clknet_1_0__leaf_net421),
    .C_N(net416),
    .D_N(net424),
    .X(net425));
 sky130_fd_sc_hd__buf_1 c431 (.A(net946),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 c432 (.A(net785),
    .X(net427));
 sky130_fd_sc_hd__and2_1 c433 (.A(net420),
    .B(net427),
    .X(net428));
 sky130_fd_sc_hd__and2_0 c434 (.A(net428),
    .B(net426),
    .X(net429));
 sky130_fd_sc_hd__and3_1 c435 (.A(net424),
    .B(net429),
    .C(net427),
    .X(net430));
 sky130_fd_sc_hd__a2111o_1 c436 (.A1(net429),
    .A2(clknet_1_0__leaf_net419),
    .B1(net428),
    .C1(clknet_1_0__leaf_net413),
    .X(net431));
 sky130_fd_sc_hd__and2_0 c437 (.A(net428),
    .B(net899),
    .X(net432));
 sky130_fd_sc_hd__or4bb_1 c438 (.A(net432),
    .B(net428),
    .C_N(net899),
    .D_N(clknet_1_0__leaf_net922),
    .X(net433));
 sky130_fd_sc_hd__or4bb_1 c439 (.A(net289),
    .B(net427),
    .C_N(net432),
    .D_N(net429),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 c44 (.A(net43),
    .X(net21));
 sky130_fd_sc_hd__and2_0 c440 (.A(net423),
    .B(net303),
    .X(net435));
 sky130_fd_sc_hd__and2_0 c441 (.A(net435),
    .B(net316),
    .X(net436));
 sky130_fd_sc_hd__buf_1 c442 (.A(clknet_1_0__leaf_net901),
    .X(net437));
 sky130_fd_sc_hd__and2_1 c443 (.A(net436),
    .B(net303),
    .X(net438));
 sky130_fd_sc_hd__buf_1 c444 (.A(clknet_1_1__leaf_net901),
    .X(net439));
 sky130_fd_sc_hd__and2_0 c445 (.A(clknet_1_0__leaf_net439),
    .B(net435),
    .X(net440));
 sky130_fd_sc_hd__and2_0 c446 (.A(net435),
    .B(clknet_1_0__leaf_net440),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 c447 (.A(net821),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 c448 (.A(net887),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 c449 (.A(net824),
    .X(net444));
 sky130_fd_sc_hd__dlymetal6s2s_1 c45 (.A(net21),
    .X(net22));
 sky130_fd_sc_hd__and2_0 c450 (.A(net443),
    .B(clknet_1_1__leaf_net439),
    .X(net445));
 sky130_fd_sc_hd__and2_0 c451 (.A(clknet_1_0__leaf_net445),
    .B(clknet_1_0__leaf_net439),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 c452 (.A(net828),
    .X(net447));
 sky130_fd_sc_hd__and2_0 c453 (.A(net446),
    .B(net444),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 c454 (.A(net833),
    .X(net449));
 sky130_fd_sc_hd__and2_0 c455 (.A(net444),
    .B(net449),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 c456 (.A(net824),
    .X(net451));
 sky130_fd_sc_hd__and2_0 c457 (.A(net442),
    .B(clknet_1_1__leaf_net445),
    .X(net452));
 sky130_fd_sc_hd__and2_0 c458 (.A(net450),
    .B(net451),
    .X(net453));
 sky130_fd_sc_hd__and2_0 c459 (.A(net453),
    .B(net451),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 c46 (.X(net768));
 sky130_fd_sc_hd__clkbuf_1 c460 (.A(net791),
    .X(net455));
 sky130_fd_sc_hd__mux4_1 c461 (.A0(net455),
    .A1(net452),
    .A2(clknet_1_0__leaf_net445),
    .A3(clknet_1_1__leaf_net448),
    .S0(clknet_1_1__leaf_net439),
    .S1(net316),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 c462 (.A(net334),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 c463 (.A(net447),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 c464 (.A(net457),
    .X(net459));
 sky130_fd_sc_hd__buf_1 c465 (.A(clknet_1_1__leaf_net901),
    .X(net460));
 sky130_fd_sc_hd__buf_1 c466 (.A(net735),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 c467 (.A(net735),
    .X(net462));
 sky130_fd_sc_hd__buf_1 c468 (.A(net820),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 c469 (.A(net1025),
    .X(net464));
 sky130_fd_sc_hd__buf_2 c47 (.A(net768),
    .X(net24));
 sky130_fd_sc_hd__buf_1 c470 (.A(net463),
    .X(net465));
 sky130_fd_sc_hd__and2_0 c471 (.A(net464),
    .B(net465),
    .X(net466));
 sky130_fd_sc_hd__and2_0 c472 (.A(net457),
    .B(net465),
    .X(net467));
 sky130_fd_sc_hd__and2_0 c473 (.A(net460),
    .B(net465),
    .X(net468));
 sky130_fd_sc_hd__or4bb_1 c474 (.A(net461),
    .B(net463),
    .C_N(net465),
    .D_N(net1053),
    .X(net469));
 sky130_fd_sc_hd__and2_1 c475 (.A(net465),
    .B(net466),
    .X(net470));
 sky130_fd_sc_hd__buf_1 c476 (.A(net1049),
    .X(net471));
 sky130_fd_sc_hd__buf_2 c477 (.A(net1038),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_1 c478 (.A(net838),
    .X(net473));
 sky130_fd_sc_hd__and2_0 c479 (.A(net322),
    .B(net472),
    .X(net474));
 sky130_fd_sc_hd__and2_0 c48 (.A(net23),
    .B(net21),
    .X(net25));
 sky130_fd_sc_hd__a2111o_1 c480 (.A1(net459),
    .A2(net470),
    .B1(net472),
    .C1(net471),
    .D1(net469),
    .X(net475));
 sky130_fd_sc_hd__sdfbbn_1 c481 (.CLK_N(clknet_4_12_0_clk),
    .D(net474),
    .RESET_B(net469),
    .SCD(net472),
    .SCE(net470),
    .SET_B(net471),
    .Q(net477),
    .Q_N(net476));
 sky130_fd_sc_hd__or4bb_1 c482 (.A(net477),
    .B(net470),
    .C_N(net471),
    .D_N(net461),
    .X(net478));
 sky130_fd_sc_hd__mux4_1 c483 (.A0(net476),
    .A1(net473),
    .A2(net470),
    .A3(net459),
    .S0(net472),
    .S1(net1066),
    .X(net479));
 sky130_fd_sc_hd__buf_1 c484 (.A(net358),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 c485 (.A(net480),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 c486 (.A(net909),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 c487 (.A(net363),
    .X(net483));
 sky130_fd_sc_hd__buf_1 c488 (.A(net358),
    .X(net484));
 sky130_fd_sc_hd__and2_1 c489 (.A(net484),
    .B(net483),
    .X(net986));
 sky130_fd_sc_hd__and2_1 c49 (.A(net21),
    .B(net20),
    .X(net26));
 sky130_fd_sc_hd__and2_0 c490 (.A(net480),
    .B(net484),
    .X(net485));
 sky130_fd_sc_hd__and3_1 c491 (.A(net482),
    .B(net485),
    .C(net484),
    .X(net486));
 sky130_fd_sc_hd__and2_1 c492 (.A(net483),
    .B(net484),
    .X(net487));
 sky130_fd_sc_hd__and2_0 c493 (.A(net481),
    .B(net483),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 c494 (.A(net890),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 c495 (.A(net890),
    .X(net490));
 sky130_fd_sc_hd__buf_1 c496 (.X(net491));
 sky130_fd_sc_hd__and2_1 c497 (.A(net489),
    .B(net491),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 c498 (.A(net814),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 c499 (.A(net782),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 c50 (.A(net780),
    .X(net27));
 sky130_fd_sc_hd__and3_1 c500 (.A(net485),
    .B(net493),
    .C(net490),
    .X(net495));
 sky130_fd_sc_hd__and2_0 c501 (.A(net491),
    .B(net494),
    .X(net496));
 sky130_fd_sc_hd__and3_1 c502 (.A(net496),
    .B(net494),
    .C(net492),
    .X(net497));
 sky130_fd_sc_hd__or4bb_1 c503 (.A(net497),
    .B(net492),
    .C_N(net495),
    .D_N(net491),
    .X(net498));
 sky130_fd_sc_hd__and3_1 c504 (.A(net480),
    .B(net489),
    .C(net890),
    .X(net499));
 sky130_fd_sc_hd__sdfxbp_1 c505 (.CLK(clknet_4_14_0_clk),
    .D(net489),
    .SCD(net495),
    .SCE(net499),
    .Q(net501),
    .Q_N(net500));
 sky130_fd_sc_hd__and2_0 c509 (.A(net388),
    .B(net500),
    .X(net502));
 sky130_fd_sc_hd__buf_1 c51 (.A(net801),
    .X(net28));
 sky130_fd_sc_hd__and2_0 c510 (.A(net502),
    .B(net1072),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 c511 (.A(net502),
    .X(net504));
 sky130_fd_sc_hd__buf_1 c512 (.A(net732),
    .X(net505));
 sky130_fd_sc_hd__and2_1 c513 (.A(net504),
    .B(net505),
    .X(net982));
 sky130_fd_sc_hd__and2_1 c514 (.A(net505),
    .B(net504),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_1 c515 (.A(net732),
    .X(net507));
 sky130_fd_sc_hd__dlymetal6s2s_1 c516 (.A(net797),
    .X(net987));
 sky130_fd_sc_hd__and3_1 c517 (.A(net507),
    .B(net987),
    .C(net500),
    .X(net508));
 sky130_fd_sc_hd__and2_1 c518 (.A(net508),
    .B(net987),
    .X(net984));
 sky130_fd_sc_hd__and2_1 c519 (.A(net503),
    .B(net505),
    .X(net509));
 sky130_fd_sc_hd__and2_0 c52 (.A(net28),
    .B(net24),
    .X(net29));
 sky130_fd_sc_hd__and2_0 c520 (.A(net502),
    .B(net388),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_1 c521 (.A(net1058),
    .X(net511));
 sky130_fd_sc_hd__and2_1 c522 (.A(net501),
    .B(net894),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 c523 (.A(net777),
    .X(net981));
 sky130_fd_sc_hd__sdfbbp_1 c524 (.CLK(clknet_4_14_0_clk),
    .D(net511),
    .RESET_B(net512),
    .SCD(net984),
    .SCE(net987),
    .SET_B(net982),
    .Q(net983),
    .Q_N(net988));
 sky130_fd_sc_hd__clkbuf_1 c525 (.A(net927),
    .X(net513));
 sky130_fd_sc_hd__and2_0 c526 (.A(net512),
    .B(net513),
    .X(net985));
 sky130_fd_sc_hd__a2111o_1 c527 (.A1(net367),
    .A2(net513),
    .B1(net987),
    .C1(net501),
    .D1(net503),
    .X(net989));
 sky130_fd_sc_hd__buf_1 c528 (.A(clknet_1_1__leaf_net922),
    .X(net514));
 sky130_fd_sc_hd__buf_1 c529 (.A(clknet_1_0__leaf_net514),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 c53 (.A(net773),
    .X(net30));
 sky130_fd_sc_hd__and2_0 c530 (.A(clknet_1_1__leaf_net515),
    .B(clknet_1_0__leaf_net514),
    .X(net516));
 sky130_fd_sc_hd__and2_0 c531 (.A(clknet_1_0__leaf_net515),
    .B(clknet_1_1__leaf_net514),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_1 c532 (.A(net743),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 c533 (.A(net742),
    .X(net519));
 sky130_fd_sc_hd__and2_0 c534 (.A(net518),
    .B(net252),
    .X(net520));
 sky130_fd_sc_hd__and2_1 c535 (.A(net520),
    .B(net518),
    .X(net521));
 sky130_fd_sc_hd__buf_1 c536 (.A(net790),
    .X(net522));
 sky130_fd_sc_hd__buf_1 c537 (.A(clknet_1_1__leaf_net514),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_1 c538 (.A(net775),
    .X(net524));
 sky130_fd_sc_hd__and2_0 c539 (.A(net524),
    .B(clknet_1_1__leaf_net523),
    .X(net525));
 sky130_fd_sc_hd__and2_1 c54 (.A(net27),
    .B(net29),
    .X(net31));
 sky130_fd_sc_hd__sdfxtp_1 c540 (.CLK(clknet_4_5_0_clk),
    .D(clknet_1_1__leaf_net525),
    .SCD(net522),
    .SCE(clknet_1_1__leaf_net523),
    .Q(net526));
 sky130_fd_sc_hd__clkbuf_1 c541 (.A(net800),
    .X(net527));
 sky130_fd_sc_hd__and2_0 c542 (.A(clknet_1_0__leaf_net523),
    .B(net520),
    .X(net528));
 sky130_fd_sc_hd__or4bb_1 c543 (.A(net521),
    .B(clknet_1_0__leaf_net525),
    .C_N(clknet_1_0__leaf_net523),
    .D_N(net992),
    .X(net529));
 sky130_fd_sc_hd__buf_1 c544 (.A(net811),
    .X(net530));
 sky130_fd_sc_hd__a2111o_1 c545 (.A1(net527),
    .A2(net530),
    .B1(clknet_1_1__leaf_net525),
    .C1(net1034),
    .D1(clknet_1_1__leaf_net523),
    .X(net531));
 sky130_fd_sc_hd__a2111o_1 c546 (.A1(net530),
    .A2(net527),
    .B1(clknet_1_0__leaf_net523),
    .C1(net992),
    .D1(net870),
    .X(net532));
 sky130_fd_sc_hd__sdfsbp_1 c547 (.CLK(clknet_4_5_0_clk),
    .D(net530),
    .SCD(clknet_1_0__leaf_net528),
    .SCE(clknet_1_1__leaf_net532),
    .SET_B(net1034),
    .Q(net534),
    .Q_N(net533));
 sky130_fd_sc_hd__and2_0 c548 (.A(net534),
    .B(net870),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 c549 (.A0(net522),
    .A1(net535),
    .A2(net533),
    .A3(net530),
    .S0(net992),
    .S1(net870),
    .X(net536));
 sky130_fd_sc_hd__and2_1 c55 (.A(net31),
    .B(net29),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 c550 (.A(net519),
    .X(net537));
 sky130_fd_sc_hd__buf_1 c551 (.A(net537),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 c552 (.A(net758),
    .X(net539));
 sky130_fd_sc_hd__and2_2 c553 (.A(net526),
    .B(net539),
    .X(net540));
 sky130_fd_sc_hd__and2_0 c554 (.A(net538),
    .B(net536),
    .X(net541));
 sky130_fd_sc_hd__and2_1 c555 (.A(net540),
    .B(net539),
    .X(net542));
 sky130_fd_sc_hd__sdfxtp_1 c556 (.CLK(clknet_4_4_0_clk),
    .D(net430),
    .SCD(net538),
    .SCE(net539),
    .Q(net543));
 sky130_fd_sc_hd__and2_1 c557 (.A(net543),
    .B(net540),
    .X(net544));
 sky130_fd_sc_hd__and2_1 c558 (.A(net544),
    .B(net543),
    .X(net545));
 sky130_fd_sc_hd__buf_1 c559 (.A(net758),
    .X(net546));
 sky130_fd_sc_hd__buf_1 c56 (.A(clknet_1_0__leaf_net943),
    .X(net33));
 sky130_fd_sc_hd__and2_0 c560 (.A(net519),
    .B(net544),
    .X(net547));
 sky130_fd_sc_hd__sdfxtp_1 c561 (.CLK(clknet_4_4_0_clk),
    .D(net541),
    .SCD(net547),
    .SCE(net544),
    .Q(net548));
 sky130_fd_sc_hd__or4bb_2 c562 (.A(net1023),
    .B(net539),
    .C_N(net992),
    .D_N(net540),
    .X(net549));
 sky130_fd_sc_hd__and2_1 c563 (.A(net542),
    .B(net549),
    .X(net550));
 sky130_fd_sc_hd__dfbbn_1 c564 (.CLK_N(clknet_4_6_0_clk),
    .D(net546),
    .RESET_B(net550),
    .SET_B(net540),
    .Q(net552),
    .Q_N(net551));
 sky130_fd_sc_hd__clkbuf_1 c565 (.A(net951),
    .X(net553));
 sky130_fd_sc_hd__a2111o_1 c566 (.A1(clknet_1_0__leaf_net532),
    .A2(net542),
    .B1(net549),
    .C1(net552),
    .D1(net540),
    .X(net554));
 sky130_fd_sc_hd__and3_1 c567 (.A(net552),
    .B(net553),
    .C(net542),
    .X(net555));
 sky130_fd_sc_hd__mux4_1 c568 (.A0(net538),
    .A1(net540),
    .A2(net539),
    .A3(net546),
    .S0(net1023),
    .S1(net550),
    .X(net556));
 sky130_fd_sc_hd__and3_1 c569 (.A(net539),
    .B(net549),
    .C(net869),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 c57 (.A0(clknet_1_0__leaf_net33),
    .A1(net23),
    .A2(net22),
    .A3(net31),
    .S0(net24),
    .S1(net28),
    .X(net34));
 sky130_fd_sc_hd__mux4_1 c570 (.A0(net547),
    .A1(net557),
    .A2(net545),
    .A3(net551),
    .S0(net546),
    .S1(net540),
    .X(net558));
 sky130_fd_sc_hd__a2111o_1 c571 (.A1(net545),
    .A2(net552),
    .B1(net543),
    .C1(net869),
    .D1(clknet_1_0__leaf_net923),
    .X(net559));
 sky130_fd_sc_hd__buf_1 c572 (.A(net536),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 c573 (.A(net744),
    .X(net561));
 sky130_fd_sc_hd__dlymetal6s2s_1 c574 (.A(net744),
    .X(net562));
 sky130_fd_sc_hd__and2_0 c575 (.A(net549),
    .B(net561),
    .X(net563));
 sky130_fd_sc_hd__buf_1 c576 (.A(net816),
    .X(net564));
 sky130_fd_sc_hd__and3_1 c577 (.A(net564),
    .B(net562),
    .C(net561),
    .X(net565));
 sky130_fd_sc_hd__and2_1 c578 (.A(net565),
    .B(net561),
    .X(net566));
 sky130_fd_sc_hd__and2_2 c579 (.A(net564),
    .B(net562),
    .X(net567));
 sky130_fd_sc_hd__sdfbbn_1 c58 (.CLK_N(clknet_4_9_0_clk),
    .D(net28),
    .RESET_B(clknet_1_1__leaf_net33),
    .SCD(net32),
    .SCE(net31),
    .SET_B(net1017),
    .Q(net36),
    .Q_N(net35));
 sky130_fd_sc_hd__clkbuf_1 c580 (.A(net947),
    .X(net568));
 sky130_fd_sc_hd__and2_1 c581 (.A(net566),
    .B(net561),
    .X(net569));
 sky130_fd_sc_hd__buf_1 c582 (.A(clknet_1_1__leaf_net898),
    .X(net570));
 sky130_fd_sc_hd__and2_0 c583 (.A(net565),
    .B(net562),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 c584 (.A(net835),
    .X(net572));
 sky130_fd_sc_hd__and2_0 c585 (.A(net568),
    .B(net561),
    .X(net573));
 sky130_fd_sc_hd__and2_0 c586 (.A(net561),
    .B(clknet_1_1__leaf_net923),
    .X(net574));
 sky130_fd_sc_hd__mux4_1 c587 (.A0(clknet_1_0__leaf_net574),
    .A1(net565),
    .A2(net562),
    .A3(net571),
    .S0(net564),
    .S1(net566),
    .X(net575));
 sky130_fd_sc_hd__buf_1 c588 (.A(net810),
    .X(net576));
 sky130_fd_sc_hd__mux4_1 c589 (.A0(net570),
    .A1(clknet_1_1__leaf_net574),
    .A2(net576),
    .A3(net565),
    .S0(net566),
    .S1(net569),
    .X(net577));
 sky130_fd_sc_hd__mux4_1 c59 (.A0(net30),
    .A1(net26),
    .A2(net31),
    .A3(net24),
    .S0(net28),
    .S1(net1017),
    .X(net37));
 sky130_fd_sc_hd__and2_0 c590 (.A(net571),
    .B(clknet_1_1__leaf_net924),
    .X(net578));
 sky130_fd_sc_hd__and2_0 c591 (.A(net576),
    .B(clknet_1_0__leaf_net924),
    .X(net579));
 sky130_fd_sc_hd__a2111o_1 c592 (.A1(net575),
    .A2(net569),
    .B1(net576),
    .C1(net562),
    .D1(net992),
    .X(net580));
 sky130_fd_sc_hd__mux4_1 c593 (.A0(net576),
    .A1(net564),
    .A2(net562),
    .A3(clknet_1_0__leaf_net898),
    .S0(clknet_1_0__leaf_net901),
    .S1(clknet_1_0__leaf_net924),
    .X(net581));
 sky130_fd_sc_hd__and2_0 c594 (.A(net572),
    .B(net472),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 c595 (.A(net471),
    .X(net583));
 sky130_fd_sc_hd__and2_1 c596 (.A(net582),
    .B(net471),
    .X(net584));
 sky130_fd_sc_hd__and2_0 c597 (.A(net579),
    .B(net584),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_1 c598 (.A(net769),
    .X(net586));
 sky130_fd_sc_hd__and2_0 c599 (.A(net582),
    .B(net471),
    .X(net587));
 sky130_fd_sc_hd__and3_1 c60 (.A(net29),
    .B(net36),
    .C(clknet_1_0__leaf_net33),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 c600 (.A(net583),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_1 c601 (.A(net769),
    .X(net589));
 sky130_fd_sc_hd__and2_0 c602 (.A(net472),
    .B(net588),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 c603 (.A(net772),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 c604 (.A(net772),
    .X(net592));
 sky130_fd_sc_hd__and2_2 c605 (.A(net588),
    .B(net582),
    .X(net593));
 sky130_fd_sc_hd__and3_1 c606 (.A(net473),
    .B(net587),
    .C(net593),
    .X(net594));
 sky130_fd_sc_hd__dfbbn_1 c607 (.CLK_N(clknet_4_13_0_clk),
    .D(net589),
    .RESET_B(net593),
    .SET_B(net914),
    .Q(net596),
    .Q_N(net595));
 sky130_fd_sc_hd__dfbbp_1 c608 (.CLK(clknet_4_13_0_clk),
    .D(net586),
    .RESET_B(net584),
    .SET_B(net593),
    .Q(net598),
    .Q_N(net597));
 sky130_fd_sc_hd__and3_1 c609 (.A(net589),
    .B(net593),
    .C(net1042),
    .X(net599));
 sky130_fd_sc_hd__and3_1 c61 (.A(net38),
    .B(net31),
    .C(net915),
    .X(net39));
 sky130_fd_sc_hd__and3_1 c610 (.A(net592),
    .B(net593),
    .C(net1030),
    .X(net600));
 sky130_fd_sc_hd__or4bb_1 c611 (.A(net591),
    .B(net598),
    .C_N(net593),
    .D_N(net1030),
    .X(net601));
 sky130_fd_sc_hd__and3_1 c612 (.A(net588),
    .B(net909),
    .C(net914),
    .X(net602));
 sky130_fd_sc_hd__sdfxbp_1 c613 (.CLK(clknet_4_13_0_clk),
    .D(net598),
    .SCD(net593),
    .SCE(net1075),
    .Q(net604),
    .Q_N(net603));
 sky130_fd_sc_hd__sdfbbn_1 c614 (.CLK_N(clknet_4_13_0_clk),
    .D(net604),
    .RESET_B(net592),
    .SCD(net593),
    .SCE(net597),
    .SET_B(net909),
    .Q(net606),
    .Q_N(net605));
 sky130_fd_sc_hd__sdfbbn_1 c615 (.CLK_N(clknet_4_13_0_clk),
    .D(net602),
    .RESET_B(net593),
    .SCD(net1063),
    .SCE(net603),
    .SET_B(net567),
    .Q(net608),
    .Q_N(net607));
 sky130_fd_sc_hd__and2_1 c616 (.A(net608),
    .B(net501),
    .X(net609));
 sky130_fd_sc_hd__and2_1 c617 (.A(net609),
    .B(net607),
    .X(net610));
 sky130_fd_sc_hd__and2_1 c618 (.A(net610),
    .B(net605),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 c619 (.A(net896),
    .X(net612));
 sky130_fd_sc_hd__and3_1 c62 (.A(net31),
    .B(net903),
    .C(net915),
    .X(net40));
 sky130_fd_sc_hd__and2_0 c620 (.A(net612),
    .B(net605),
    .X(net613));
 sky130_fd_sc_hd__and2_1 c621 (.A(net613),
    .B(net612),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_1 c622 (.A(net895),
    .X(net615));
 sky130_fd_sc_hd__and2_0 c623 (.A(net613),
    .B(net615),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 c624 (.A(net789),
    .X(net617));
 sky130_fd_sc_hd__and2_1 c625 (.A(net614),
    .B(net609),
    .X(net618));
 sky130_fd_sc_hd__and2_1 c626 (.A(net615),
    .B(net613),
    .X(net991));
 sky130_fd_sc_hd__and2_0 c627 (.A(net501),
    .B(net991),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_1 c628 (.A(net809),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 c629 (.A(net808),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_1 c63 (.A(net1021),
    .X(net41));
 sky130_fd_sc_hd__and2_0 c630 (.A(net621),
    .B(net596),
    .X(net622));
 sky130_fd_sc_hd__and2_1 c631 (.A(net620),
    .B(net612),
    .X(net623));
 sky130_fd_sc_hd__and2_0 c632 (.A(net622),
    .B(net623),
    .X(net624));
 sky130_fd_sc_hd__buf_1 c633 (.A(net912),
    .X(net625));
 sky130_fd_sc_hd__and3_1 c634 (.A(net617),
    .B(net625),
    .C(net620),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_1 c635 (.A(net881),
    .X(net626));
 sky130_fd_sc_hd__mux4_1 c636 (.A0(net619),
    .A1(net625),
    .A2(net622),
    .A3(net623),
    .S0(net621),
    .S1(clknet_1_1__leaf_net923),
    .X(net627));
 sky130_fd_sc_hd__mux4_2 c637 (.A0(net624),
    .A1(net626),
    .A2(net990),
    .A3(net623),
    .S0(net625),
    .S1(net896),
    .X(net980));
 sky130_fd_sc_hd__and3_1 c64 (.A(net32),
    .B(net41),
    .C(net40),
    .X(net42));
 sky130_fd_sc_hd__buf_1 c65 (.A(net20),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 c66 (.A(net902),
    .X(net44));
 sky130_fd_sc_hd__buf_1 c660 (.A(net992),
    .X(net628));
 sky130_fd_sc_hd__and2_2 c661 (.A(net628),
    .B(net992),
    .X(net629));
 sky130_fd_sc_hd__and3_1 c662 (.A(net629),
    .B(net628),
    .C(net536),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_1 c663 (.A(net748),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 c664 (.A(net748),
    .X(net632));
 sky130_fd_sc_hd__and2_1 c665 (.A(net1057),
    .B(net629),
    .X(net633));
 sky130_fd_sc_hd__and2_0 c666 (.A(net632),
    .B(net631),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 c667 (.A(net776),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 c668 (.A(net813),
    .X(net636));
 sky130_fd_sc_hd__and2_1 c669 (.A(net634),
    .B(net636),
    .X(net637));
 sky130_fd_sc_hd__buf_1 c67 (.A(net44),
    .X(net45));
 sky130_fd_sc_hd__sdfxbp_1 c670 (.CLK(clknet_4_5_0_clk),
    .D(net630),
    .SCD(net637),
    .SCE(net629),
    .Q(net639),
    .Q_N(net638));
 sky130_fd_sc_hd__clkbuf_1 c671 (.A(net836),
    .X(net640));
 sky130_fd_sc_hd__and2_1 c672 (.A(net639),
    .B(net632),
    .X(net641));
 sky130_fd_sc_hd__and2_2 c673 (.A(net641),
    .B(net631),
    .X(net642));
 sky130_fd_sc_hd__and3_1 c674 (.A(net635),
    .B(net639),
    .C(net642),
    .X(net643));
 sky130_fd_sc_hd__buf_1 c675 (.A(net953),
    .X(net644));
 sky130_fd_sc_hd__mux4_1 c676 (.A0(net643),
    .A1(net638),
    .A2(net630),
    .A3(net644),
    .S0(net628),
    .S1(net629),
    .X(net645));
 sky130_fd_sc_hd__or4bb_1 c677 (.A(net640),
    .B(net644),
    .C_N(net642),
    .D_N(net629),
    .X(net646));
 sky130_fd_sc_hd__mux4_1 c678 (.A0(net644),
    .A1(net638),
    .A2(net642),
    .A3(net629),
    .S0(net646),
    .S1(net1037),
    .X(net647));
 sky130_fd_sc_hd__mux4_1 c679 (.A0(net646),
    .A1(net642),
    .A2(net629),
    .A3(net643),
    .S1(net926),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_2 c68 (.A(net45),
    .X(net46));
 sky130_fd_sc_hd__sdfbbp_1 c680 (.CLK(clknet_4_7_0_clk),
    .D(net636),
    .RESET_B(net630),
    .SCD(net642),
    .SCE(net868),
    .SET_B(net925),
    .Q(net650),
    .Q_N(net649));
 sky130_fd_sc_hd__and3_1 c681 (.A(net649),
    .B(net634),
    .C(net868),
    .X(net651));
 sky130_fd_sc_hd__and2_0 c682 (.A(net650),
    .B(clknet_1_0__leaf_net923),
    .X(net652));
 sky130_fd_sc_hd__sdfxtp_1 c683 (.CLK(clknet_4_7_0_clk),
    .D(net298),
    .SCD(net651),
    .SCE(net992),
    .Q(net653));
 sky130_fd_sc_hd__buf_1 c684 (.A(net939),
    .X(net654));
 sky130_fd_sc_hd__and2_0 c685 (.A(clknet_1_0__leaf_net652),
    .B(clknet_1_0__leaf_net923),
    .X(net655));
 sky130_fd_sc_hd__and2_0 c686 (.A(net651),
    .B(net654),
    .X(net656));
 sky130_fd_sc_hd__and2_0 c687 (.A(clknet_1_0__leaf_net655),
    .B(clknet_1_0__leaf_net652),
    .X(net657));
 sky130_fd_sc_hd__buf_1 c688 (.A(net764),
    .X(net658));
 sky130_fd_sc_hd__sdfxtp_1 c689 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net655),
    .SCD(clknet_1_1__leaf_net657),
    .SCE(net658),
    .Q(net659));
 sky130_fd_sc_hd__buf_1 c69 (.A(net731),
    .X(net47));
 sky130_fd_sc_hd__and3_1 c690 (.A(net659),
    .B(clknet_1_1__leaf_net652),
    .C(clknet_1_1__leaf_net655),
    .X(net660));
 sky130_fd_sc_hd__and2_1 c691 (.A(net654),
    .B(net659),
    .X(net661));
 sky130_fd_sc_hd__and3_1 c692 (.A(net656),
    .B(clknet_1_0__leaf_net660),
    .C(clknet_1_1__leaf_net652),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_1 c693 (.A(net763),
    .X(net663));
 sky130_fd_sc_hd__sdfsbp_1 c694 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net657),
    .SCD(net1079),
    .SCE(clknet_1_0__leaf_net652),
    .SET_B(clknet_1_0__leaf_net923),
    .Q(net665),
    .Q_N(net664));
 sky130_fd_sc_hd__and3_1 c695 (.A(net654),
    .B(net665),
    .C(clknet_1_1__leaf_net655),
    .X(net666));
 sky130_fd_sc_hd__buf_1 c696 (.A(net784),
    .X(net667));
 sky130_fd_sc_hd__and3_1 c697 (.A(net663),
    .B(net659),
    .C(net667),
    .X(net668));
 sky130_fd_sc_hd__and3_1 c698 (.A(net658),
    .B(net654),
    .C(net668),
    .X(net669));
 sky130_fd_sc_hd__and3_1 c699 (.A(net668),
    .B(net667),
    .C(clknet_1_0__leaf_net666),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 c70 (.A(net731),
    .X(net48));
 sky130_fd_sc_hd__a2111o_1 c700 (.A1(net653),
    .A2(net661),
    .B1(net667),
    .C1(clknet_1_1__leaf_net652),
    .D1(net875),
    .X(net671));
 sky130_fd_sc_hd__or4bb_1 c701 (.A(net664),
    .B(net654),
    .C_N(clknet_1_1__leaf_net666),
    .D_N(net876),
    .X(net672));
 sky130_fd_sc_hd__and3_1 c702 (.A(net665),
    .B(net671),
    .C(clknet_1_1__leaf_net655),
    .X(net673));
 sky130_fd_sc_hd__mux4_1 c703 (.A0(net673),
    .A1(clknet_1_1__leaf_net660),
    .A2(net668),
    .A3(clknet_1_1__leaf_net655),
    .S0(clknet_1_1__leaf_net652),
    .X(net674));
 sky130_fd_sc_hd__dlymetal6s2s_1 c704 (.A(net573),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 c705 (.A(net888),
    .X(net676));
 sky130_fd_sc_hd__and2_1 c706 (.A(net669),
    .B(net567),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 c707 (.A(net888),
    .X(net678));
 sky130_fd_sc_hd__and2_0 c708 (.A(net676),
    .B(net661),
    .X(net679));
 sky130_fd_sc_hd__and2_0 c709 (.A(net661),
    .B(net910),
    .X(net680));
 sky130_fd_sc_hd__and2_0 c71 (.A(net47),
    .B(net45),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 c710 (.A(net567),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_2 c711 (.A(net1039),
    .X(net682));
 sky130_fd_sc_hd__and2_0 c712 (.A(net679),
    .B(net682),
    .X(net683));
 sky130_fd_sc_hd__and2_0 c713 (.A(net678),
    .B(net675),
    .X(net684));
 sky130_fd_sc_hd__and2_0 c714 (.A(net680),
    .B(net682),
    .X(net685));
 sky130_fd_sc_hd__buf_1 c715 (.A(clknet_1_0__leaf_net898),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_1 c716 (.A(net828),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_1 c717 (.A(net887),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 c718 (.A(net813),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_1 c719 (.A(net787),
    .X(net690));
 sky130_fd_sc_hd__and2_1 c72 (.A(net44),
    .B(net1061),
    .X(net50));
 sky130_fd_sc_hd__and2_1 c720 (.A(net689),
    .B(net682),
    .X(net691));
 sky130_fd_sc_hd__and3_1 c721 (.A(net690),
    .B(net682),
    .C(net691),
    .X(net692));
 sky130_fd_sc_hd__buf_1 c722 (.A(net783),
    .X(net693));
 sky130_fd_sc_hd__and3_1 c723 (.A(net692),
    .B(net688),
    .C(net693),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 c724 (.A(net954),
    .X(net695));
 sky130_fd_sc_hd__and2_0 c725 (.A(net695),
    .B(net693),
    .X(net696));
 sky130_fd_sc_hd__buf_1 c726 (.A(net596),
    .X(net697));
 sky130_fd_sc_hd__dlymetal6s2s_1 c727 (.A(net606),
    .X(net698));
 sky130_fd_sc_hd__and2_0 c728 (.A(net697),
    .B(net698),
    .X(net699));
 sky130_fd_sc_hd__buf_1 c729 (.A(net698),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 c73 (.A(net826),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 c730 (.A(net698),
    .X(net701));
 sky130_fd_sc_hd__and2_1 c731 (.A(net699),
    .B(net698),
    .X(net702));
 sky130_fd_sc_hd__and2_1 c732 (.A(net701),
    .B(net682),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_1 c733 (.A(net765),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_1 c734 (.A(net765),
    .X(net705));
 sky130_fd_sc_hd__and2_0 c735 (.A(net696),
    .B(net700),
    .X(net706));
 sky130_fd_sc_hd__sdfxtp_1 c736 (.CLK(clknet_4_13_0_clk),
    .D(net706),
    .SCD(net702),
    .SCE(net698),
    .Q(net707));
 sky130_fd_sc_hd__and2_0 c737 (.A(net682),
    .B(net704),
    .X(net708));
 sky130_fd_sc_hd__dfbbn_1 c738 (.CLK_N(clknet_4_7_0_clk),
    .D(net702),
    .RESET_B(net700),
    .SET_B(net682),
    .Q(net710),
    .Q_N(net709));
 sky130_fd_sc_hd__dfbbn_1 c739 (.CLK_N(clknet_4_13_0_clk),
    .D(net708),
    .RESET_B(net703),
    .SET_B(net1062),
    .Q(net712),
    .Q_N(net711));
 sky130_fd_sc_hd__clkbuf_1 c74 (.A(net795),
    .X(net52));
 sky130_fd_sc_hd__and3_1 c740 (.A(net710),
    .B(net708),
    .C(net707),
    .X(net713));
 sky130_fd_sc_hd__and3_1 c741 (.A(net705),
    .B(net710),
    .C(net712),
    .X(net714));
 sky130_fd_sc_hd__and3_1 c742 (.A(net697),
    .B(net714),
    .C(net709),
    .X(net715));
 sky130_fd_sc_hd__a2111o_1 c743 (.A1(net714),
    .A2(net710),
    .B1(net707),
    .C1(net661),
    .D1(net698),
    .X(net716));
 sky130_fd_sc_hd__and3_1 c744 (.A(net713),
    .B(net715),
    .C(net716),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 c745 (.A(net882),
    .X(net718));
 sky130_fd_sc_hd__or4bb_1 c746 (.A(net712),
    .B(net707),
    .C_N(net716),
    .D_N(net709),
    .X(net719));
 sky130_fd_sc_hd__mux4_1 c747 (.A0(net704),
    .A1(net719),
    .A2(net714),
    .A3(net716),
    .S0(net595),
    .S1(net697),
    .X(net720));
 sky130_fd_sc_hd__buf_1 c748 (.X(net750));
 sky130_fd_sc_hd__clkbuf_2 c749 (.A(net751),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 c75 (.A(net807),
    .X(net53));
 sky130_fd_sc_hd__sdfstp_1 c750 (.CLK(clknet_4_15_0_clk),
    .D(net990),
    .SCD(net722),
    .SCE(net980),
    .SET_B(net472),
    .Q(net723));
 sky130_fd_sc_hd__sdfstp_1 c751 (.CLK(clknet_4_15_0_clk),
    .D(net722),
    .SCD(net1070),
    .SCE(net980),
    .SET_B(net721),
    .Q(net724));
 sky130_fd_sc_hd__a2111o_1 c752 (.A1(net723),
    .A2(net990),
    .B1(net724),
    .C1(net722),
    .D1(net882),
    .X(net725));
 sky130_fd_sc_hd__and3_1 c753 (.A(net724),
    .B(net725),
    .C(net722),
    .X(net726));
 sky130_fd_sc_hd__sdfbbn_1 c754 (.CLK_N(clknet_4_15_0_clk),
    .D(net675),
    .RESET_B(net726),
    .SCD(net724),
    .SCE(net725),
    .SET_B(net722),
    .Q(net728),
    .Q_N(net727));
 sky130_fd_sc_hd__a2111o_1 c755 (.A1(net728),
    .A2(net723),
    .B1(net726),
    .C1(net722),
    .D1(net724),
    .X(net729));
 sky130_fd_sc_hd__mux4_1 c756 (.A0(net726),
    .A1(net725),
    .A2(net727),
    .A3(net722),
    .S0(net724),
    .S1(net913),
    .X(net730));
 sky130_fd_sc_hd__and2_1 c76 (.A(net48),
    .B(net45),
    .X(net54));
 sky130_fd_sc_hd__and2_1 c77 (.A(net50),
    .B(net51),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 c78 (.A(net812),
    .X(net56));
 sky130_fd_sc_hd__sdfrbp_1 c79 (.CLK(clknet_4_8_0_clk),
    .D(net46),
    .RESET_B(net54),
    .SCD(net43),
    .SCE(net55),
    .Q(net58),
    .Q_N(net57));
 sky130_fd_sc_hd__clkbuf_1 c80 (.A(net931),
    .X(net59));
 sky130_fd_sc_hd__sdfbbp_1 c81 (.CLK(clknet_4_10_0_clk),
    .D(net52),
    .RESET_B(net55),
    .SCD(net45),
    .SCE(net56),
    .SET_B(net47),
    .Q(net61),
    .Q_N(net60));
 sky130_fd_sc_hd__and3_1 c82 (.A(net53),
    .B(net59),
    .C(net60),
    .X(net62));
 sky130_fd_sc_hd__and2_1 c83 (.A(net61),
    .B(net56),
    .X(net63));
 sky130_fd_sc_hd__a2111o_1 c84 (.A1(net59),
    .A2(net62),
    .B1(net63),
    .C1(net60),
    .D1(net55),
    .X(net64));
 sky130_fd_sc_hd__a2111o_1 c85 (.A1(net51),
    .A2(net63),
    .B1(net56),
    .C1(net1048),
    .D1(net891),
    .X(net65));
 sky130_fd_sc_hd__or4bb_1 c86 (.A(net49),
    .B(net65),
    .C_N(net1082),
    .D_N(net1048),
    .X(net66));
 sky130_fd_sc_hd__or4bb_1 c87 (.A(net47),
    .B(net62),
    .C_N(net63),
    .D_N(net891),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 c88 (.A(net24),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 c89 (.A(net68),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 c90 (.A(net68),
    .X(net70));
 sky130_fd_sc_hd__and2_0 c91 (.A(net58),
    .B(net69),
    .X(net71));
 sky130_fd_sc_hd__and2_1 c92 (.A(net43),
    .B(net68),
    .X(net72));
 sky130_fd_sc_hd__and2_0 c93 (.A(net70),
    .B(net72),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 c94 (.X(net747));
 sky130_fd_sc_hd__and2_0 c95 (.A(net69),
    .B(net72),
    .X(net75));
 sky130_fd_sc_hd__and2_0 c96 (.A(net74),
    .B(net72),
    .X(net76));
 sky130_fd_sc_hd__buf_1 c97 (.A(net747),
    .X(net77));
 sky130_fd_sc_hd__and2_1 c98 (.A(net77),
    .B(net74),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 c99 (.A(net779),
    .X(net79));
 sky130_fd_sc_hd__buf_1 merge757 (.A(net1058),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 merge758 (.A(net802),
    .X(net732));
 sky130_fd_sc_hd__dfbbp_1 merge759 (.CLK(clknet_4_0_0_clk),
    .D(net250),
    .RESET_B(net127),
    .SET_B(net253),
    .Q(net734),
    .Q_N(net733));
 sky130_fd_sc_hd__clkbuf_1 merge760 (.A(net1025),
    .X(net735));
 sky130_fd_sc_hd__or4bb_1 merge761 (.A(net578),
    .B(net661),
    .C_N(net581),
    .D_N(net677),
    .X(net736));
 sky130_fd_sc_hd__sdfxbp_1 merge762 (.CLK(clknet_4_1_0_clk),
    .D(clknet_1_0__leaf_net415),
    .SCD(net285),
    .SCE(clknet_1_0__leaf_net413),
    .Q(net738),
    .Q_N(net737));
 sky130_fd_sc_hd__sdfbbn_1 merge763 (.CLK_N(clknet_4_5_0_clk),
    .D(net397),
    .RESET_B(net399),
    .SCD(net391),
    .SCE(net392),
    .SET_B(net390),
    .Q(net740),
    .Q_N(net739));
 sky130_fd_sc_hd__or4bb_1 merge764 (.A(net114),
    .B(net119),
    .C_N(net121),
    .D_N(net124),
    .X(net741));
 sky130_fd_sc_hd__sdfxbp_1 merge765 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net516),
    .SCD(clknet_1_1__leaf_net514),
    .SCE(net517),
    .Q(net743),
    .Q_N(net742));
 sky130_fd_sc_hd__buf_1 merge766 (.A(net940),
    .X(net744));
 sky130_fd_sc_hd__buf_1 merge767 (.A(clknet_1_1__leaf_net794),
    .X(net745));
 sky130_fd_sc_hd__or4bb_1 merge768 (.A(net434),
    .B(net316),
    .C_N(net437),
    .D_N(net430),
    .X(net746));
 sky130_fd_sc_hd__sdfstp_1 merge769 (.CLK(clknet_4_8_0_clk),
    .D(net71),
    .SCD(net72),
    .SCE(net73),
    .Q(net747));
 sky130_fd_sc_hd__clkbuf_1 merge770 (.A(net787),
    .X(net748));
 sky130_fd_sc_hd__sdfxtp_1 merge771 (.CLK(clknet_4_10_0_clk),
    .D(net109),
    .SCD(net231),
    .SCE(net210),
    .Q(net749));
 sky130_fd_sc_hd__sedfxbp_1 merge772 (.CLK(clknet_4_15_0_clk),
    .DE(net980),
    .SCD(net718),
    .SCE(net500),
    .Q(net751),
    .Q_N(net750));
 sky130_fd_sc_hd__or4bb_1 merge773 (.A(net609),
    .B(net986),
    .C_N(net611),
    .D_N(net500),
    .X(net752));
 sky130_fd_sc_hd__sedfxbp_1 merge774 (.CLK(clknet_4_14_0_clk),
    .D(net357),
    .DE(net365),
    .SCD(net369),
    .Q(net368),
    .Q_N(net753));
 sky130_fd_sc_hd__buf_1 merge775 (.A(net803),
    .X(net755));
 sky130_fd_sc_hd__sedfxtp_1 merge776 (.CLK(clknet_4_2_0_clk),
    .D(net5),
    .DE(net3),
    .SCD(net0),
    .SCE(net2),
    .Q(net756));
 sky130_fd_sc_hd__sedfxtp_2 merge777 (.CLK(clknet_4_8_0_clk),
    .D(net75),
    .DE(net90),
    .SCD(net95),
    .Q(net92));
 sky130_fd_sc_hd__clkbuf_1 merge778 (.A(net934),
    .X(net758));
 sky130_fd_sc_hd__buf_1 merge779 (.A(clknet_1_1__leaf_net944),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 merge780 (.A(net780),
    .X(net760));
 sky130_fd_sc_hd__sedfxtp_1 merge781 (.CLK(clknet_4_9_0_clk),
    .D(net39),
    .DE(net144),
    .SCD(net162),
    .SCE(clknet_1_1__leaf_net164),
    .Q(net761));
 sky130_fd_sc_hd__and3_1 merge782 (.A(net488),
    .B(net485),
    .C(net486),
    .X(net762));
 sky130_fd_sc_hd__sdfrbp_1 merge783 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net657),
    .RESET_B(clknet_1_1__leaf_net652),
    .SCD(clknet_1_0__leaf_net660),
    .SCE(clknet_1_0__leaf_net655),
    .Q(net764),
    .Q_N(net763));
 sky130_fd_sc_hd__clkbuf_1 merge784 (.A(net932),
    .X(net765));
 sky130_fd_sc_hd__sdfrbp_1 merge785 (.CLK(clknet_4_11_0_clk),
    .D(net189),
    .RESET_B(net202),
    .SCD(net207),
    .SCE(net205),
    .Q(net767),
    .Q_N(net766));
 sky130_fd_sc_hd__sdfxtp_1 merge786 (.CLK(clknet_4_8_0_clk),
    .D(net43),
    .SCD(net22),
    .Q(net768));
 sky130_fd_sc_hd__clkbuf_1 merge787 (.A(net952),
    .X(net769));
 sky130_fd_sc_hd__sdfrtn_1 merge788 (.CLK_N(clknet_4_11_0_clk),
    .D(net198),
    .RESET_B(clknet_1_0__leaf_net321),
    .SCE(net323),
    .Q(net322));
 sky130_fd_sc_hd__sdfrtp_1 merge789 (.CLK(clknet_4_3_0_clk),
    .D(net145),
    .RESET_B(net144),
    .SCD(net154),
    .SCE(net277),
    .Q(net771));
 sky130_fd_sc_hd__clkbuf_1 merge790 (.A(net913),
    .X(net772));
 sky130_fd_sc_hd__sdfrtp_1 merge791 (.CLK(clknet_4_12_0_clk),
    .D(clknet_1_0__leaf_net138),
    .RESET_B(net1051),
    .SCD(net26),
    .SCE(net22),
    .Q(net773));
 sky130_fd_sc_hd__sdfrtp_1 merge792 (.CLK(clknet_4_12_0_clk),
    .D(net141),
    .RESET_B(net1051),
    .SCE(net142),
    .Q(net143));
 sky130_fd_sc_hd__sdfsbp_1 merge793 (.CLK(clknet_4_5_0_clk),
    .D(net628),
    .SCD(net630),
    .SCE(net399),
    .SET_B(clknet_1_1__leaf_net523),
    .Q(net776),
    .Q_N(net775));
 sky130_fd_sc_hd__sdfsbp_1 merge794 (.CLK(clknet_4_15_0_clk),
    .D(net468),
    .SCD(net459),
    .SCE(net506),
    .SET_B(net509),
    .Q(net778),
    .Q_N(net777));
 sky130_fd_sc_hd__sdfstp_1 merge795 (.CLK(clknet_4_8_0_clk),
    .D(net63),
    .SCD(net71),
    .SCE(net76),
    .SET_B(net86),
    .Q(net779));
 sky130_fd_sc_hd__buf_1 merge796 (.A(net942),
    .X(net780));
 sky130_fd_sc_hd__sdfstp_1 merge797 (.CLK(clknet_4_3_0_clk),
    .D(net281),
    .SCD(net144),
    .SCE(net299),
    .SET_B(clknet_1_0__leaf_net302),
    .Q(net781));
 sky130_fd_sc_hd__sdfstp_1 merge798 (.CLK(clknet_4_11_0_clk),
    .D(net184),
    .SCD(net185),
    .SCE(net487),
    .SET_B(net492),
    .Q(net782));
 sky130_fd_sc_hd__sedfxbp_1 merge799 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_0__leaf_net666),
    .DE(net658),
    .SCD(net685),
    .SCE(net691),
    .Q(net784),
    .Q_N(net783));
 sky130_fd_sc_hd__sedfxbp_1 merge800 (.CLK(clknet_4_1_0_clk),
    .D(net146),
    .DE(net144),
    .SCD(clknet_1_1__leaf_net419),
    .SCE(net426),
    .Q(net786),
    .Q_N(net785));
 sky130_fd_sc_hd__sedfxtp_1 merge801 (.CLK(clknet_4_7_0_clk),
    .D(net630),
    .DE(net629),
    .SCD(net687),
    .SCE(net677),
    .Q(net787));
 sky130_fd_sc_hd__or4bb_1 merge802 (.A(clknet_1_0__leaf_net686),
    .B(net677),
    .C_N(clknet_1_0__leaf_net441),
    .D_N(clknet_1_1__leaf_net440),
    .X(net788));
 sky130_fd_sc_hd__sedfxtp_1 merge803 (.CLK(clknet_4_15_0_clk),
    .D(net329),
    .DE(net323),
    .SCD(net611),
    .SCE(net614),
    .Q(net789));
 sky130_fd_sc_hd__sedfxtp_1 merge804 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_1__leaf_net413),
    .DE(clknet_1_1__leaf_net421),
    .SCD(clknet_1_1__leaf_net516),
    .SCE(net521),
    .Q(net790));
 sky130_fd_sc_hd__sdfrbp_1 merge805 (.CLK(clknet_4_3_0_clk),
    .D(net137),
    .RESET_B(net144),
    .SCD(net438),
    .SCE(net454),
    .Q(net792),
    .Q_N(net791));
 sky130_fd_sc_hd__a2111o_1 merge806 (.A1(net114),
    .A2(net113),
    .B1(net112),
    .C1(net118),
    .D1(net964),
    .X(net793));
 sky130_fd_sc_hd__buf_1 merge807 (.A(clknet_1_0__leaf_net944),
    .X(net794));
 sky130_fd_sc_hd__sdfrbp_1 merge808 (.CLK(clknet_4_10_0_clk),
    .D(net201),
    .RESET_B(net209),
    .SCD(net48),
    .SCE(net46),
    .Q(net796),
    .Q_N(net795));
 sky130_fd_sc_hd__sdfrtn_1 merge809 (.CLK_N(clknet_4_14_0_clk),
    .D(net355),
    .RESET_B(net353),
    .SCD(net505),
    .SCE(net506),
    .Q(net797));
 sky130_fd_sc_hd__sdfxtp_1 merge810 (.CLK(clknet_4_10_0_clk),
    .D(net237),
    .SCD(net231),
    .SCE(net1045),
    .Q(net798));
 sky130_fd_sc_hd__sdfrtp_1 merge811 (.CLK(clknet_4_12_0_clk),
    .D(net459),
    .RESET_B(net461),
    .SCD(net323),
    .SCE(net463),
    .Q(net799));
 sky130_fd_sc_hd__sdfrtp_1 merge812 (.CLK(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net525),
    .RESET_B(clknet_1_0__leaf_net523),
    .SCD(clknet_1_1__leaf_net415),
    .SCE(net422),
    .Q(net800));
 sky130_fd_sc_hd__sdfrtp_1 merge813 (.CLK(clknet_4_9_0_clk),
    .D(net25),
    .RESET_B(net23),
    .SCD(net173),
    .SCE(net172),
    .Q(net801));
 sky130_fd_sc_hd__sdfbbp_1 merge814 (.CLK(clknet_4_14_0_clk),
    .D(net347),
    .RESET_B(net345),
    .SCD(net504),
    .SCE(net986),
    .SET_B(net982),
    .Q(net803),
    .Q_N(net802));
 sky130_fd_sc_hd__dfbbn_1 merge815 (.CLK_N(clknet_4_4_0_clk),
    .D(clknet_1_0__leaf_net415),
    .RESET_B(net418),
    .SET_B(clknet_1_0__leaf_net421),
    .Q(net805),
    .Q_N(net804));
 sky130_fd_sc_hd__sdfsbp_1 merge816 (.CLK(clknet_4_10_0_clk),
    .D(net49),
    .SCD(net50),
    .SCE(net193),
    .SET_B(net191),
    .Q(net807),
    .Q_N(net806));
 sky130_fd_sc_hd__sdfbbn_1 merge817 (.CLK_N(clknet_4_15_0_clk),
    .D(net616),
    .RESET_B(net619),
    .SCD(net617),
    .SCE(net618),
    .SET_B(net991),
    .Q(net809),
    .Q_N(net808));
 sky130_fd_sc_hd__sdfsbp_1 merge818 (.CLK(clknet_4_7_0_clk),
    .D(clknet_1_1__leaf_net528),
    .SCD(net522),
    .SCE(net569),
    .SET_B(net567),
    .Q(net811),
    .Q_N(net810));
 sky130_fd_sc_hd__sdfstp_1 merge819 (.CLK(clknet_4_10_0_clk),
    .D(net99),
    .SCD(net98),
    .SCE(net54),
    .SET_B(net50),
    .Q(net812));
 sky130_fd_sc_hd__sdfstp_1 merge820 (.CLK(clknet_4_7_0_clk),
    .D(net633),
    .SCD(net635),
    .SCE(net683),
    .SET_B(net682),
    .Q(net813));
 sky130_fd_sc_hd__sdfbbn_1 merge821 (.CLK_N(clknet_4_14_0_clk),
    .D(net486),
    .RESET_B(net1052),
    .SCD(net986),
    .SCE(net488),
    .Q(net491),
    .Q_N(net814));
 sky130_fd_sc_hd__sdfstp_1 merge822 (.CLK(clknet_4_6_0_clk),
    .D(net681),
    .SCD(net677),
    .SCE(net563),
    .SET_B(net1040),
    .Q(net816));
 sky130_fd_sc_hd__or4bb_1 merge823 (.A(net300),
    .B(clknet_1_0__leaf_net301),
    .C_N(net335),
    .D_N(net330),
    .X(net817));
 sky130_fd_sc_hd__sedfxbp_1 merge824 (.CLK(clknet_4_11_0_clk),
    .D(clknet_1_1__leaf_net321),
    .DE(net329),
    .SCD(net181),
    .SCE(net184),
    .Q(net819),
    .Q_N(net818));
 sky130_fd_sc_hd__sedfxbp_1 merge825 (.CLK(clknet_4_6_0_clk),
    .D(clknet_1_1__leaf_net439),
    .DE(net438),
    .SCD(net458),
    .SCE(net459),
    .Q(net821),
    .Q_N(net820));
 sky130_fd_sc_hd__sdfbbp_1 merge826 (.CLK(clknet_4_2_0_clk),
    .D(net205),
    .RESET_B(net212),
    .SCD(net119),
    .SCE(net122),
    .SET_B(net127),
    .Q(net823),
    .Q_N(net822));
 sky130_fd_sc_hd__sedfxtp_1 merge827 (.CLK(clknet_4_6_0_clk),
    .D(net449),
    .DE(clknet_1_0__leaf_net448),
    .SCD(clknet_1_0__leaf_net440),
    .SCE(net438),
    .Q(net824));
 sky130_fd_sc_hd__sedfxtp_1 merge828 (.CLK(clknet_4_10_0_clk),
    .D(net97),
    .DE(net95),
    .SCD(net101),
    .SCE(net98),
    .Q(net825));
 sky130_fd_sc_hd__sdfbbn_1 merge829 (.CLK_N(clknet_4_10_0_clk),
    .D(net98),
    .RESET_B(net99),
    .SCD(net45),
    .SCE(net46),
    .SET_B(net50),
    .Q(net827),
    .Q_N(net826));
 sky130_fd_sc_hd__sedfxtp_1 merge830 (.CLK(clknet_4_6_0_clk),
    .D(net436),
    .DE(clknet_1_1__leaf_net441),
    .SCD(net677),
    .SCE(clknet_1_1__leaf_net686),
    .Q(net828));
 sky130_fd_sc_hd__mux4_1 merge831 (.A0(net324),
    .A1(net325),
    .A2(net323),
    .A3(net510),
    .S0(net512),
    .S1(net509),
    .X(net829));
 sky130_fd_sc_hd__mux4_1 merge832 (.A0(net241),
    .A1(net239),
    .A2(net185),
    .A3(net183),
    .S0(net187),
    .S1(net879),
    .X(net830));
 sky130_fd_sc_hd__mux4_1 merge833 (.A0(net243),
    .A1(net231),
    .A2(net241),
    .A3(net55),
    .S0(net53),
    .S1(net57),
    .X(net831));
 sky130_fd_sc_hd__sdfbbn_1 merge834 (.CLK_N(clknet_4_3_0_clk),
    .D(clknet_1_0__leaf_net448),
    .RESET_B(net444),
    .SCD(clknet_1_1__leaf_net302),
    .SCE(net303),
    .SET_B(net300),
    .Q(net833),
    .Q_N(net832));
 sky130_fd_sc_hd__or4bb_1 merge835 (.A(net562),
    .B(net560),
    .C_N(net684),
    .D_N(net682),
    .X(net834));
 sky130_fd_sc_hd__sdfrbp_1 merge836 (.CLK(clknet_4_7_0_clk),
    .D(net637),
    .RESET_B(net633),
    .SCD(net569),
    .SCE(net566),
    .Q(net836),
    .Q_N(net835));
 sky130_fd_sc_hd__mux4_1 merge837 (.A0(net394),
    .A1(net392),
    .A2(net391),
    .A3(net700),
    .S0(net703),
    .S1(net702),
    .X(net837));
 sky130_fd_sc_hd__sdfbbp_1 merge838 (.CLK(clknet_4_13_0_clk),
    .D(net462),
    .RESET_B(net458),
    .SCD(net470),
    .SCE(net467),
    .SET_B(net465),
    .Q(net839),
    .Q_N(net838));
 sky130_fd_sc_hd__mux4_1 merge839 (.A0(net341),
    .A1(clknet_1_0__leaf_net321),
    .A2(net128),
    .A3(net126),
    .S0(net113),
    .S1(net907),
    .X(net840));
 sky130_fd_sc_hd__mux4_1 merge840 (.A0(net433),
    .A1(net545),
    .A2(net539),
    .A3(net393),
    .S0(net397),
    .S1(net389),
    .X(net841));
 sky130_fd_sc_hd__mux4_1 merge841 (.A0(net316),
    .A1(net335),
    .A2(net326),
    .A3(net380),
    .S0(net373),
    .S1(net379),
    .X(net842));
 sky130_fd_sc_hd__mux4_1 merge842 (.A0(net313),
    .A1(net316),
    .A2(clknet_1_0__leaf_net310),
    .A3(net124),
    .S0(net121),
    .S1(net127),
    .X(net843));
 sky130_fd_sc_hd__mux4_1 merge843 (.A0(clknet_1_0__leaf_net652),
    .A1(net653),
    .A2(net434),
    .A3(net130),
    .S0(net132),
    .S1(net117),
    .X(net844));
 sky130_fd_sc_hd__mux4_1 merge844 (.A0(net144),
    .A1(net282),
    .A2(net281),
    .A3(net560),
    .S0(net908),
    .S1(clknet_1_0__leaf_net923),
    .X(net845));
 sky130_fd_sc_hd__mux4_1 merge845 (.A0(net35),
    .A1(net46),
    .A2(net47),
    .A3(net509),
    .S0(net984),
    .S1(net1072),
    .X(net846));
 sky130_fd_sc_hd__mux4_1 merge846 (.A0(net179),
    .A1(net24),
    .A2(net25),
    .A3(net330),
    .S0(net323),
    .S1(net907),
    .X(net847));
 sky130_fd_sc_hd__mux4_1 merge847 (.A0(net22),
    .A1(net32),
    .A2(net31),
    .A3(net368),
    .S0(net384),
    .S1(net382),
    .X(net848));
 sky130_fd_sc_hd__mux4_1 merge848 (.A0(net716),
    .A1(net717),
    .A2(net711),
    .A3(net623),
    .S0(net610),
    .S1(net611),
    .X(net849));
 sky130_fd_sc_hd__mux4_1 merge849 (.A0(net134),
    .A1(net127),
    .A2(clknet_1_0__leaf_net135),
    .A3(net300),
    .S0(net285),
    .S1(clknet_1_0__leaf_net302),
    .X(net850));
 sky130_fd_sc_hd__mux4_1 merge850 (.A0(net127),
    .A1(net253),
    .A2(net252),
    .A3(net126),
    .S0(net254),
    .S1(net250),
    .X(net851));
 sky130_fd_sc_hd__mux4_1 merge851 (.A0(net560),
    .A1(net566),
    .A2(net561),
    .A3(net416),
    .S0(net423),
    .S1(clknet_1_1__leaf_net421),
    .X(net852));
 sky130_fd_sc_hd__mux4_1 merge852 (.A0(net208),
    .A1(net218),
    .A2(net216),
    .A3(net379),
    .S0(net382),
    .S1(net373),
    .X(net853));
 sky130_fd_sc_hd__mux4_1 merge853 (.A0(net550),
    .A1(net551),
    .A2(net549),
    .A3(net308),
    .S0(clknet_1_1__leaf_net307),
    .S1(net305),
    .X(net854));
 sky130_fd_sc_hd__sdfbbn_1 merge854 (.CLK_N(clknet_4_9_0_clk),
    .D(clknet_1_0__leaf_net164),
    .RESET_B(net159),
    .SCD(clknet_1_0__leaf_net157),
    .SCE(net166),
    .SET_B(net163),
    .Q(net856),
    .Q_N(net855));
 sky130_fd_sc_hd__mux4_1 merge855 (.A0(clknet_1_1__leaf_net310),
    .A1(net300),
    .A2(clknet_1_1__leaf_net307),
    .A3(net555),
    .S0(net584),
    .S1(clknet_1_0__leaf_net585),
    .X(net857));
 sky130_fd_sc_hd__mux4_1 merge856 (.A0(net642),
    .A1(net643),
    .A2(net641),
    .A3(net259),
    .S0(net252),
    .S1(net997),
    .X(net858));
 sky130_fd_sc_hd__mux4_1 merge857 (.A0(net142),
    .A1(net146),
    .A2(net144),
    .A3(net694),
    .S0(net693),
    .S1(net691),
    .X(net859));
 sky130_fd_sc_hd__mux4_1 merge858 (.A0(net326),
    .A1(net323),
    .A2(net322),
    .A3(net377),
    .S0(net367),
    .S1(net379),
    .X(net860));
 sky130_fd_sc_hd__mux4_1 merge859 (.A0(net349),
    .A1(net354),
    .A2(net357),
    .A3(net40),
    .S0(net32),
    .S1(net35),
    .X(net861));
 sky130_fd_sc_hd__mux4_1 merge860 (.A0(clknet_1_1__leaf_net585),
    .A1(net587),
    .A2(net590),
    .A3(net350),
    .S0(net623),
    .S1(net618),
    .X(net862));
 sky130_fd_sc_hd__mux4_1 merge861 (.A0(net392),
    .A1(net391),
    .A2(net394),
    .A3(net389),
    .S0(net397),
    .S1(net399),
    .X(net863));
 sky130_fd_sc_hd__dfrbp_1 merge862 (.CLK(clknet_4_12_0_clk),
    .D(net360),
    .RESET_B(net361),
    .Q(net865),
    .Q_N(net864));
 sky130_fd_sc_hd__dfrbp_1 merge863 (.CLK(clknet_4_8_0_clk),
    .D(net221),
    .RESET_B(net225),
    .Q(net867),
    .Q_N(net866));
 sky130_fd_sc_hd__dfrtn_1 merge864 (.CLK_N(clknet_4_5_0_clk),
    .D(net647),
    .Q(net868));
 sky130_fd_sc_hd__dfrtp_1 merge865 (.CLK(clknet_4_6_0_clk),
    .D(net554),
    .RESET_B(net1024),
    .Q(net869));
 sky130_fd_sc_hd__dfrtp_1 merge866 (.CLK(clknet_4_5_0_clk),
    .D(net529),
    .RESET_B(net531),
    .Q(net870));
 sky130_fd_sc_hd__dfrtp_1 merge867 (.CLK(clknet_4_12_0_clk),
    .D(net152),
    .RESET_B(net1028),
    .Q(net871));
 sky130_fd_sc_hd__dfsbp_1 merge868 (.CLK(clknet_4_2_0_clk),
    .D(net167),
    .SET_B(net176),
    .Q(net873),
    .Q_N(net872));
 sky130_fd_sc_hd__and2_0 merge869 (.A(net730),
    .B(net729),
    .X(net874));
 sky130_fd_sc_hd__dfsbp_1 merge870 (.CLK(clknet_4_7_0_clk),
    .D(net662),
    .SET_B(net670),
    .Q(net876),
    .Q_N(net875));
 sky130_fd_sc_hd__and2_0 merge871 (.A(net600),
    .B(net1031),
    .X(net877));
 sky130_fd_sc_hd__dfstp_1 merge872 (.CLK(clknet_4_4_0_clk),
    .D(net402),
    .SET_B(net403),
    .Q(net878));
 sky130_fd_sc_hd__dfstp_1 merge873 (.CLK(clknet_4_10_0_clk),
    .D(net242),
    .SET_B(net1036),
    .Q(net879));
 sky130_fd_sc_hd__dfstp_1 merge874 (.CLK(clknet_4_0_0_clk),
    .D(net741),
    .SET_B(net793),
    .Q(net880));
 sky130_fd_sc_hd__dlrbn_1 merge875 (.D(net720),
    .GATE_N(clknet_4_15_0_clk),
    .RESET_B(net849),
    .Q(net882),
    .Q_N(net881));
 sky130_fd_sc_hd__dlrbn_1 merge876 (.D(net262),
    .GATE_N(clknet_4_1_0_clk),
    .RESET_B(net270),
    .Q(net884),
    .Q_N(net883));
 sky130_fd_sc_hd__dlrbp_1 merge877 (.D(net192),
    .GATE(clknet_4_11_0_clk),
    .RESET_B(net200),
    .Q(net886),
    .Q_N(net885));
 sky130_fd_sc_hd__dlrbp_1 merge878 (.D(net736),
    .GATE(clknet_4_6_0_clk),
    .RESET_B(net788),
    .Q(net888),
    .Q_N(net887));
 sky130_fd_sc_hd__dlrtn_1 merge879 (.D(net319),
    .GATE_N(clknet_4_9_0_clk),
    .RESET_B(net817),
    .Q(net889));
 sky130_fd_sc_hd__dlrtn_1 merge880 (.D(net498),
    .GATE_N(clknet_4_14_0_clk),
    .RESET_B(net762),
    .Q(net890));
 sky130_fd_sc_hd__dlrtn_1 merge881 (.D(net64),
    .GATE_N(clknet_4_10_0_clk),
    .RESET_B(net66),
    .Q(net891));
 sky130_fd_sc_hd__dlrtp_1 merge882 (.D(net287),
    .GATE(clknet_4_3_0_clk),
    .RESET_B(net297),
    .Q(net892));
 sky130_fd_sc_hd__dlrtp_1 merge883 (.D(net107),
    .GATE(clknet_4_10_0_clk),
    .RESET_B(net103),
    .Q(net893));
 sky130_fd_sc_hd__dlrtp_1 merge884 (.D(net374),
    .GATE(clknet_4_14_0_clk),
    .RESET_B(net376),
    .Q(net894));
 sky130_fd_sc_hd__edfxbp_1 merge885 (.CLK(clknet_4_15_0_clk),
    .D(net627),
    .DE(net752),
    .Q(net896),
    .Q_N(net895));
 sky130_fd_sc_hd__edfxtp_1 merge886 (.CLK(clknet_4_2_0_clk),
    .D(net14),
    .DE(net18),
    .Q(net897));
 sky130_fd_sc_hd__sdlclkp_1 merge887 (.CLK(clknet_4_6_0_clk),
    .GATE(net580),
    .SCE(net834),
    .GCLK(net898));
 sky130_fd_sc_hd__sdlclkp_2 merge888 (.CLK(clknet_4_4_0_clk),
    .GATE(net425),
    .GCLK(net431));
 sky130_fd_sc_hd__and2_1 merge889 (.A(net339),
    .B(net340),
    .X(net900));
 sky130_fd_sc_hd__sdlclkp_4 merge890 (.CLK(clknet_4_6_0_clk),
    .GATE(net456),
    .SCE(net746),
    .GCLK(net901));
 sky130_fd_sc_hd__dfrbp_1 merge891 (.CLK(clknet_4_9_0_clk),
    .D(net37),
    .RESET_B(net1022),
    .Q(net903),
    .Q_N(net902));
 sky130_fd_sc_hd__dfrbp_1 merge892 (.CLK(clknet_4_13_0_clk),
    .D(net475),
    .RESET_B(net478),
    .Q(net905),
    .Q_N(net904));
 sky130_fd_sc_hd__dfrtn_1 merge893 (.CLK_N(clknet_4_8_0_clk),
    .D(net89),
    .RESET_B(net84),
    .Q(net906));
 sky130_fd_sc_hd__dfrtp_4 merge894 (.CLK(clknet_4_8_0_clk),
    .D(net900),
    .RESET_B(net16),
    .Q(net907));
 sky130_fd_sc_hd__dfrtp_1 merge895 (.CLK(clknet_4_1_0_clk),
    .D(net272),
    .RESET_B(net559),
    .Q(net908));
 sky130_fd_sc_hd__dfrtp_1 merge896 (.CLK(clknet_4_15_0_clk),
    .D(net479),
    .RESET_B(net877),
    .Q(net909));
 sky130_fd_sc_hd__dfsbp_1 merge897 (.CLK(clknet_4_7_0_clk),
    .D(net672),
    .Q(net674),
    .Q_N(net910));
 sky130_fd_sc_hd__dfsbp_1 merge898 (.CLK(clknet_4_15_0_clk),
    .D(net874),
    .SET_B(net862),
    .Q(net913),
    .Q_N(net912));
 sky130_fd_sc_hd__dfstp_1 merge899 (.CLK(clknet_4_13_0_clk),
    .D(net594),
    .SET_B(net599),
    .Q(net914));
 sky130_fd_sc_hd__dfxbp_1 s900 (.CLK(clknet_4_9_0_clk),
    .D(net34),
    .Q(net916),
    .Q_N(net915));
 sky130_fd_sc_hd__dfxbp_1 s901 (.CLK(clknet_4_10_0_clk),
    .D(net108),
    .Q(net918),
    .Q_N(net917));
 sky130_fd_sc_hd__dfxtp_1 s902 (.CLK(clknet_4_10_0_clk),
    .D(net111),
    .Q(net919));
 sky130_fd_sc_hd__dfxtp_1 s903 (.CLK(clknet_4_11_0_clk),
    .D(net249),
    .Q(net920));
 sky130_fd_sc_hd__dfxtp_1 s904 (.CLK(clknet_4_5_0_clk),
    .D(net408),
    .Q(net921));
 sky130_fd_sc_hd__dlclkp_1 s905 (.CLK(clknet_4_4_0_clk),
    .GATE(net412),
    .GCLK(net922));
 sky130_fd_sc_hd__dlclkp_2 s906 (.CLK(clknet_4_6_0_clk),
    .GATE(net558),
    .GCLK(net923));
 sky130_fd_sc_hd__dlclkp_4 s907 (.CLK(clknet_4_6_0_clk),
    .GATE(net577),
    .GCLK(net924));
 sky130_fd_sc_hd__dlxbn_1 s908 (.D(net645),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net926),
    .Q_N(net925));
 sky130_fd_sc_hd__dlxbn_1 s909 (.D(net829),
    .GATE_N(clknet_4_14_0_clk),
    .Q(net928),
    .Q_N(net927));
 sky130_fd_sc_hd__dlxbp_1 s910 (.D(net830),
    .GATE(clknet_4_11_0_clk),
    .Q(net930),
    .Q_N(net929));
 sky130_fd_sc_hd__dlxtn_1 s911 (.D(net831),
    .GATE_N(clknet_4_10_0_clk),
    .Q(net931));
 sky130_fd_sc_hd__dlxtn_1 s912 (.D(net837),
    .GATE_N(clknet_4_5_0_clk),
    .Q(net932));
 sky130_fd_sc_hd__dlxtn_4 s913 (.D(net840),
    .GATE_N(clknet_4_2_0_clk),
    .Q(net933));
 sky130_fd_sc_hd__dlxtp_1 s914 (.D(net841),
    .GATE(clknet_4_4_0_clk),
    .Q(net934));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s915 (.D(net842),
    .SLEEP_B(clknet_4_11_0_clk),
    .Q(net935));
 sky130_fd_sc_hd__dfxbp_1 s916 (.CLK(clknet_4_2_0_clk),
    .D(net843),
    .Q(net937),
    .Q_N(net936));
 sky130_fd_sc_hd__dfxbp_1 s917 (.CLK(clknet_4_3_0_clk),
    .D(net844),
    .Q(net939),
    .Q_N(net938));
 sky130_fd_sc_hd__dfxtp_1 s918 (.CLK(clknet_4_1_0_clk),
    .D(net845),
    .Q(net940));
 sky130_fd_sc_hd__dfxtp_1 s919 (.CLK(clknet_4_11_0_clk),
    .D(net846),
    .Q(net941));
 sky130_fd_sc_hd__dfxtp_1 s920 (.CLK(clknet_4_9_0_clk),
    .D(net847),
    .Q(net942));
 sky130_fd_sc_hd__dlclkp_1 s921 (.CLK(clknet_4_9_0_clk),
    .GATE(net848),
    .GCLK(net943));
 sky130_fd_sc_hd__dlclkp_2 s922 (.CLK(clknet_4_12_0_clk),
    .GATE(net850),
    .GCLK(net944));
 sky130_fd_sc_hd__dlclkp_4 s923 (.CLK(clknet_4_0_0_clk),
    .GATE(net851),
    .GCLK(net945));
 sky130_fd_sc_hd__dlxbn_1 s924 (.D(net852),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net947),
    .Q_N(net946));
 sky130_fd_sc_hd__dlxbn_1 s925 (.D(net853),
    .GATE_N(clknet_4_9_0_clk),
    .Q(net949),
    .Q_N(net948));
 sky130_fd_sc_hd__dlxbp_1 s926 (.D(net854),
    .GATE(clknet_4_3_0_clk),
    .Q(net951),
    .Q_N(net950));
 sky130_fd_sc_hd__dlxtn_1 s927 (.D(net857),
    .GATE_N(clknet_4_12_0_clk),
    .Q(net952));
 sky130_fd_sc_hd__dlxtn_1 s928 (.D(net858),
    .GATE_N(clknet_4_1_0_clk),
    .Q(net953));
 sky130_fd_sc_hd__dlxtn_1 s929 (.D(net859),
    .GATE_N(clknet_4_6_0_clk),
    .Q(net954));
 sky130_fd_sc_hd__dlxtp_1 s930 (.D(net860),
    .GATE(clknet_4_11_0_clk),
    .Q(net955));
 sky130_fd_sc_hd__lpflow_inputisolatch_1 s931 (.D(net861),
    .SLEEP_B(clknet_4_12_0_clk),
    .Q(net956));
 sky130_fd_sc_hd__dfxbp_1 s932 (.CLK(clknet_4_5_0_clk),
    .D(net863),
    .Q(net958),
    .Q_N(net957));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(in0),
    .X(net648));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in10),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in11),
    .X(net911));
 sky130_fd_sc_hd__buf_1 input5 (.A(in12),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in13),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(in14),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in15),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(in16),
    .X(net963));
 sky130_fd_sc_hd__buf_1 input10 (.A(in17),
    .X(net964));
 sky130_fd_sc_hd__buf_1 input11 (.A(in18),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in19),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(in2),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(in20),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(in21),
    .X(net969));
 sky130_fd_sc_hd__buf_1 input16 (.A(in22),
    .X(net970));
 sky130_fd_sc_hd__buf_1 input17 (.A(in23),
    .X(net971));
 sky130_fd_sc_hd__buf_1 input18 (.A(in24),
    .X(net972));
 sky130_fd_sc_hd__buf_1 input19 (.A(in3),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(in4),
    .X(net974));
 sky130_fd_sc_hd__buf_1 input21 (.A(in5),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in6),
    .X(net976));
 sky130_fd_sc_hd__buf_1 input23 (.A(in7),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in8),
    .X(net978));
 sky130_fd_sc_hd__buf_1 input25 (.A(in9),
    .X(net979));
 sky130_fd_sc_hd__buf_2 output26 (.A(net980),
    .X(out15));
 sky130_fd_sc_hd__buf_2 output27 (.A(net981),
    .X(out16));
 sky130_fd_sc_hd__buf_2 output28 (.A(net982),
    .X(out19));
 sky130_fd_sc_hd__buf_2 output29 (.A(net983),
    .X(out2));
 sky130_fd_sc_hd__buf_2 output30 (.A(net984),
    .X(out21));
 sky130_fd_sc_hd__buf_2 output31 (.A(net985),
    .X(out22));
 sky130_fd_sc_hd__buf_2 output32 (.A(net986),
    .X(out23));
 sky130_fd_sc_hd__buf_2 output33 (.A(net987),
    .X(out24));
 sky130_fd_sc_hd__buf_2 output34 (.A(net988),
    .X(out3));
 sky130_fd_sc_hd__buf_2 output35 (.A(net989),
    .X(out4));
 sky130_fd_sc_hd__buf_2 output36 (.A(net990),
    .X(out6));
 sky130_fd_sc_hd__buf_2 output37 (.A(net991),
    .X(out9));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net526),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net945 (.A(net945),
    .X(clknet_0_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_0__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net945 (.A(clknet_0_net945),
    .X(clknet_1_1__leaf_net945));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net260 (.A(net260),
    .X(clknet_0_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_0__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net260 (.A(clknet_0_net260),
    .X(clknet_1_1__leaf_net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net255 (.A(net255),
    .X(clknet_0_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_0__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net255 (.A(clknet_0_net255),
    .X(clknet_1_1__leaf_net255));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net944 (.A(net944),
    .X(clknet_0_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_0__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net944 (.A(clknet_0_net944),
    .X(clknet_1_1__leaf_net944));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net794 (.A(net794),
    .X(clknet_0_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_0__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net794 (.A(clknet_0_net794),
    .X(clknet_1_1__leaf_net794));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net745 (.A(net745),
    .X(clknet_0_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net745 (.A(clknet_0_net745),
    .X(clknet_1_0__leaf_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net745 (.A(clknet_0_net745),
    .X(clknet_1_1__leaf_net745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net302 (.A(net302),
    .X(clknet_0_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_0__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net302 (.A(clknet_0_net302),
    .X(clknet_1_1__leaf_net302));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net301 (.A(net301),
    .X(clknet_0_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_0__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net301 (.A(clknet_0_net301),
    .X(clknet_1_1__leaf_net301));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net321 (.A(net321),
    .X(clknet_0_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net321 (.A(clknet_0_net321),
    .X(clknet_1_1__leaf_net321));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net307 (.A(net307),
    .X(clknet_0_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_0__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net307 (.A(clknet_0_net307),
    .X(clknet_1_1__leaf_net307));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net310 (.A(net310),
    .X(clknet_0_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_0__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net310 (.A(clknet_0_net310),
    .X(clknet_1_1__leaf_net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net759 (.A(net759),
    .X(clknet_0_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_0__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net759 (.A(clknet_0_net759),
    .X(clknet_1_1__leaf_net759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net138 (.A(net138),
    .X(clknet_0_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_0__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net138 (.A(clknet_0_net138),
    .X(clknet_1_1__leaf_net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net135 (.A(net135),
    .X(clknet_0_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_0__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net135 (.A(clknet_0_net135),
    .X(clknet_1_1__leaf_net135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net157 (.A(net157),
    .X(clknet_0_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_0__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net157 (.A(clknet_0_net157),
    .X(clknet_1_1__leaf_net157));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net178 (.A(net178),
    .X(clknet_0_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_0__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net178 (.A(clknet_0_net178),
    .X(clknet_1_1__leaf_net178));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net196 (.A(net196),
    .X(clknet_0_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_0__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net196 (.A(clknet_0_net196),
    .X(clknet_1_1__leaf_net196));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net164 (.A(net164),
    .X(clknet_0_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_0__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net164 (.A(clknet_0_net164),
    .X(clknet_1_1__leaf_net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net943 (.A(net943),
    .X(clknet_0_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net943 (.A(clknet_0_net943),
    .X(clknet_1_0__leaf_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net943 (.A(clknet_0_net943),
    .X(clknet_1_1__leaf_net943));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net33 (.A(net33),
    .X(clknet_0_net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net33 (.A(clknet_0_net33),
    .X(clknet_1_0__leaf_net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net33 (.A(clknet_0_net33),
    .X(clknet_1_1__leaf_net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net924 (.A(net924),
    .X(clknet_0_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_0__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net924 (.A(clknet_0_net924),
    .X(clknet_1_1__leaf_net924));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net585 (.A(net585),
    .X(clknet_0_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_0__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net585 (.A(clknet_0_net585),
    .X(clknet_1_1__leaf_net585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net923 (.A(net923),
    .X(clknet_0_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net923 (.A(clknet_0_net923),
    .X(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net655 (.A(net655),
    .X(clknet_0_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_0__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net655 (.A(clknet_0_net655),
    .X(clknet_1_1__leaf_net655));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net666 (.A(net666),
    .X(clknet_0_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net666 (.A(clknet_0_net666),
    .X(clknet_1_0__leaf_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net666 (.A(clknet_0_net666),
    .X(clknet_1_1__leaf_net666));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net660 (.A(net660),
    .X(clknet_0_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_0__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net660 (.A(clknet_0_net660),
    .X(clknet_1_1__leaf_net660));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net657 (.A(net657),
    .X(clknet_0_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_0__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net657 (.A(clknet_0_net657),
    .X(clknet_1_1__leaf_net657));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net652 (.A(net652),
    .X(clknet_0_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net652 (.A(clknet_0_net652),
    .X(clknet_1_1__leaf_net652));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net574 (.A(net574),
    .X(clknet_0_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_0__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net574 (.A(clknet_0_net574),
    .X(clknet_1_1__leaf_net574));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net898 (.A(net898),
    .X(clknet_0_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_0__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net898 (.A(clknet_0_net898),
    .X(clknet_1_1__leaf_net898));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net686 (.A(net686),
    .X(clknet_0_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_0__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net686 (.A(clknet_0_net686),
    .X(clknet_1_1__leaf_net686));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net922 (.A(net922),
    .X(clknet_0_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_0__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net922 (.A(clknet_0_net922),
    .X(clknet_1_1__leaf_net922));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net514 (.A(net514),
    .X(clknet_0_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_0__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net514 (.A(clknet_0_net514),
    .X(clknet_1_1__leaf_net514));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net523 (.A(net523),
    .X(clknet_0_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_0__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net523 (.A(clknet_0_net523),
    .X(clknet_1_1__leaf_net523));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net532 (.A(net532),
    .X(clknet_0_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_0__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net532 (.A(clknet_0_net532),
    .X(clknet_1_1__leaf_net532));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net528 (.A(net528),
    .X(clknet_0_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_0__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net528 (.A(clknet_0_net528),
    .X(clknet_1_1__leaf_net528));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net525 (.A(net525),
    .X(clknet_0_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_0__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net525 (.A(clknet_0_net525),
    .X(clknet_1_1__leaf_net525));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net516 (.A(net516),
    .X(clknet_0_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_0__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net516 (.A(clknet_0_net516),
    .X(clknet_1_1__leaf_net516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net515 (.A(net515),
    .X(clknet_0_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_0__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net515 (.A(clknet_0_net515),
    .X(clknet_1_1__leaf_net515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net413 (.A(net413),
    .X(clknet_0_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_0__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net413 (.A(clknet_0_net413),
    .X(clknet_1_1__leaf_net413));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net421 (.A(net421),
    .X(clknet_0_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_0__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net421 (.A(clknet_0_net421),
    .X(clknet_1_1__leaf_net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net414 (.A(net414),
    .X(clknet_0_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net414 (.A(clknet_0_net414),
    .X(clknet_1_0__leaf_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net414 (.A(clknet_0_net414),
    .X(clknet_1_1__leaf_net414));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net419 (.A(net419),
    .X(clknet_0_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_0__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net419 (.A(clknet_0_net419),
    .X(clknet_1_1__leaf_net419));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net415 (.A(net415),
    .X(clknet_0_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_0__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net415 (.A(clknet_0_net415),
    .X(clknet_1_1__leaf_net415));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net901 (.A(net901),
    .X(clknet_0_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_0__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net901 (.A(clknet_0_net901),
    .X(clknet_1_1__leaf_net901));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net439 (.A(net439),
    .X(clknet_0_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_0__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net439 (.A(clknet_0_net439),
    .X(clknet_1_1__leaf_net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net448 (.A(net448),
    .X(clknet_0_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_0__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net448 (.A(clknet_0_net448),
    .X(clknet_1_1__leaf_net448));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net445 (.A(net445),
    .X(clknet_0_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_0__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net445 (.A(clknet_0_net445),
    .X(clknet_1_1__leaf_net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net440 (.A(net440),
    .X(clknet_0_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_0__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net440 (.A(clknet_0_net440),
    .X(clknet_1_1__leaf_net440));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net441 (.A(net441),
    .X(clknet_0_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_0__leaf_net441));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net441 (.A(clknet_0_net441),
    .X(clknet_1_1__leaf_net441));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer1 (.A(net998),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net264),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net994),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net253),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net253),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net1000),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net1006),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer15 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer16 (.A(net933),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net916),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net383),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net266),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net223),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net956),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net42),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net548),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net556),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net799),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net143),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net154),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net155),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net267),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net914),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net601),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net217),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net364),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net992),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net232),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net246),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net926),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net778),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net816),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net561),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net92),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net597),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net919),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net801),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net233),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net367),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net375),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net58),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net839),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net865),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net139),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net490),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net322),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net11),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net373),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net921),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net631),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net941),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net934),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net291),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net24),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net709),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net606),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net265),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net756),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net905),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net893),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net894),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net892),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net723),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net866),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net388),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net263),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net867),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net904),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net917),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net883),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net407),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net653),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net781),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net222),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net61),
    .X(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(in0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in11));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in13));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in15));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(in17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(in18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(in19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(in2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(in20));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(in21));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(in22));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(in23));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(in24));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(in3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(in4));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(in5));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(in6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(in7));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(in8));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(in9));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge806_B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_S1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_C (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c138_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c137_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c135_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c134_B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c133_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_c132_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_SCE (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c409_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c146_A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_c142_X (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_SET_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_RESET_B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_SCE (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_c147_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_DE (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_SCD (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_RESET_B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_DE (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c175_D_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c172_D1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_c164_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge857_A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge800_D (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_c308_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c204_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c197_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_Q_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_c289_C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_D (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_SCE (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c237_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_SCD (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_RESET_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_SET_B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_c224_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_RESET_B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_D (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_c230_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold69_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c88_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c59_A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c57_S0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c52_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c47_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c183_B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c181_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_c267_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c271_C (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_S0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge850_A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c534_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c410_D1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c398_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c396_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c288_B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c282_D1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_c266_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge849_S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge762_SCD (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_SCE (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c299_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c297_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_c307_X (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_SCE (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c443_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c440_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c347_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_C_N (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_D_N (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c321_B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c314_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_c312_X (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge842_A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge841_A0 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge768_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c461_S1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c441_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c329_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c328_D_N (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c327_B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_Q (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold61_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_Q (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c360_B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_C (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c337_B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c333_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_c331_X (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge858_A1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_S0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge831_A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge811_SCD (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_DE (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_SCE (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c349_S1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_c332_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_A3 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge823_D_N (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c341_B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c339_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_c462_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c382_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c358_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c348_C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c344_B (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c343_X (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_c354_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_c351_X (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge845_A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_SCE (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_SCE (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c68_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_SET_B (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c602_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c594_B (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c483_S0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c481_SCD (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c480_B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c479_B (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_c477_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge851_A0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_A3 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge835_B (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_c572_X (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_SET_B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c710_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c706_B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c615_SET_B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_c579_X (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge855_S0 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c608_RESET_B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c597_B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_c596_X (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_A0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_SCD (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c678_A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c677_C_N (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_C (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_c673_X (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge856_A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c679_A3 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c676_A0 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_c674_X (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold87_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c700_A1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_Q (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c713_B (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_c704_X (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_RESET_B (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c735_B (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_c729_X (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_S1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_D (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c736_SCD (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_c731_X (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge837_S0 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c739_RESET_B (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_c732_X (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_Q (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge846_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_SET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_c42_S1 (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_Q (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge784_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_c402_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_c161_B (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_c170_C (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_c166_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_c141_B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold42_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_X (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_SCE (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c592_D1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c562_C_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c661_B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c660_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c549_S0 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c546_C1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_c543_D_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c279_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c280_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c303_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c36_CLK_N (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge759_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge874_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s923_CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_X (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c43_CLK_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge776_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge826_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge868_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge886_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s913_GATE_N (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s916_CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_X (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c301_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c325_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge789_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge797_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge805_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge834_CLK_N (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge882_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s917_CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s926_GATE (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_X (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c540_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c547_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c670_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge763_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge793_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge864_CLK_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge866_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s904_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s908_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s912_GATE_N (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s932_CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_X (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c564_CLK_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge822_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge825_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge827_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge830_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge865_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge878_GATE (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge887_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge890_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s906_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s907_CLK (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s924_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s929_GATE_N (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_X (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c680_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c683_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c689_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c738_CLK_N (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge783_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge799_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge801_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge818_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge820_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge836_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge870_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge897_CLK (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_X (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c238_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c79_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge769_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge777_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge786_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge795_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge863_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge893_CLK_N (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge894_CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_X (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c231_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c233_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c241_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c58_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge781_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge813_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge854_CLK_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge879_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge891_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s900_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s920_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s921_CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s925_GATE_N (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_X (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c229_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c247_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c248_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c252_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c81_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge771_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge808_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge810_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge816_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge819_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge828_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge829_CLK_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge873_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge881_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge883_GATE (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s901_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s902_CLK (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s911_GATE_N (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_X (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c218_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c395_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge785_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_CLK_N (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge798_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge824_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge877_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s903_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s910_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s915_SLEEP_B (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s919_CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s930_GATE (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_X (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c367_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c380_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c385_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c387_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c390_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c505_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c524_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge774_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge809_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge814_CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge821_CLK_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge880_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge884_GATE (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_s909_GATE_N (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_X (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c750_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c751_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_c754_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge772_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge794_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge803_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge817_CLK_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge875_GATE_N (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge885_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge896_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge898_CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_X (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge788_RESET_B (.DIODE(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge839_A1 (.DIODE(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net321_X (.DIODE(clknet_1_0__leaf_net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_c571_D1 (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c682_B (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_B (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SET_B (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge844_S1 (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net923_X (.DIODE(clknet_1_0__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c586_B (.DIODE(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c636_S1 (.DIODE(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_net923_X (.DIODE(clknet_1_1__leaf_net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_c685_A (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c687_B (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_c694_SCE (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_merge843_A0 (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_net652_X (.DIODE(clknet_1_0__leaf_net652));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net979));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
